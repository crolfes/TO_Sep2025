** Created by: circuit_gen.AN2D1_1
** Cell name: AN2D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_AN2D1_1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
M_u2_M_u3 net6 a1 x_u2_net6 vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u3_M_u2 z net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u2_M_u4 x_u2_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u3_M_u3 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u2 net6 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u1 net6 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AN2D1_2
** Cell name: AN2D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_AN2D1_2 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
M_u2_M_u3 net6 a1 x_u2_net6 vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u3_M_u2 z net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u2_M_u4 x_u2_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u3_M_u3 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u2 net6 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u1 net6 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AN2D1_3
** Cell name: AN2D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_AN2D1_3 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
M_u2_M_u3 net6 a1 x_u2_net6 vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u3_M_u2 z net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u2_M_u4 x_u2_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u3_M_u3 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u2 net6 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u1 net6 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AN2D1
** Cell name: AN2D1
** Lib name: sg13g2
.SUBCKT sg13g2_AN2D1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
M_u2_M_u3 net6 a1 x_u2_net6 vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u3_M_u2 z net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u2_M_u4 x_u2_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u3_M_u3 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u2 net6 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u1 net6 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AO21D1_1
** Cell name: AO21D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_AO21D1_1 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI7 net32 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u7 net59 a1 net32 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI6 net59 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI8_M_u2 z net59 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u3 net22 a1 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI8_M_u3 z net59 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u4 net22 a2 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net22 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AO21D1_2
** Cell name: AO21D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_AO21D1_2 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI7 net32 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u7 net59 a1 net32 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI6 net59 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI8_M_u2 z net59 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u3 net22 a1 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI8_M_u3 z net59 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u4 net22 a2 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net22 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AO21D1_3
** Cell name: AO21D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_AO21D1_3 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI7 net32 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u7 net59 a1 net32 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI6 net59 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI8_M_u2 z net59 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u3 net22 a1 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI8_M_u3 z net59 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u4 net22 a2 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net22 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AO21D1
** Cell name: AO21D1
** Lib name: sg13g2
.SUBCKT sg13g2_AO21D1 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI7 net32 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u7 net59 a1 net32 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI6 net59 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI8_M_u2 z net59 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u3 net22 a1 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI8_M_u3 z net59 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u4 net22 a2 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net22 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AOI21D1_1
** Cell name: AOI21D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_AOI21D1_1 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
MI2 zn a1 net27 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI3 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u7 zn b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u4 net13 a2 zn vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net13 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u3 net13 a1 zn vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AOI21D1_2
** Cell name: AOI21D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_AOI21D1_2 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
MI2 zn a1 net27 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI3 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u7 zn b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u4 net13 a2 zn vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net13 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u3 net13 a1 zn vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AOI21D1_3
** Cell name: AOI21D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_AOI21D1_3 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
MI2 zn a1 net27 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI3 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u7 zn b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u4 net13 a2 zn vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net13 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u3 net13 a1 zn vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.AOI21D1
** Cell name: AOI21D1
** Lib name: sg13g2
.SUBCKT sg13g2_AOI21D1 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
MI2 zn a1 net27 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI3 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u7 zn b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u4 net13 a2 zn vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net13 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u3 net13 a1 zn vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ANTENNA
** Cell name: ANTENNA
** Lib name: sg13g2f
.SUBCKT sg13g2_ANTENNA i vdd vss
*.PININFO i:I vdd:B vss:B
Ddn_1 vss i dantenna m=1 w=1.485u l=970n a=1440.45f
DD0 i vdd dpantenna m=1 w=1.485u l=970n a=1440.45f
.ENDS


******* EOF

** Created by: circuit_gen.BUFFD1_1
** Cell name: BUFFD1_1
** Lib name: sg13g2
.SUBCKT sg13g2_BUFFD1_1 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u3_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u2_M_u2 net8 i vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u3_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u3 net8 i vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.BUFFD1_2
** Cell name: BUFFD1_2
** Lib name: sg13g2
.SUBCKT sg13g2_BUFFD1_2 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u3_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u2_M_u2 net8 i vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u3_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u3 net8 i vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.BUFFD1_3
** Cell name: BUFFD1_3
** Lib name: sg13g2
.SUBCKT sg13g2_BUFFD1_3 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u3_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u2_M_u2 net8 i vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u3_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u3 net8 i vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.BUFFD1
** Cell name: BUFFD1
** Lib name: sg13g2
.SUBCKT sg13g2_BUFFD1 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u3_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u2_M_u2 net8 i vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u3_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2_M_u3 net8 i vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.DFCNQD1
** Cell name: DFCNQD1
** Lib name: sg13g2
.SUBCKT sg13g2_DFCNQD1 cdn cp d q vdd vss
*.PININFO cdn:I cp:I d:I q:O vdd:B vss:B 
Mcpbn incpb cp vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07 $pos=0 $flip=0
Mcpbp incpb cp vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07 $pos=0 $flip=0
Mcpn incp incpb vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07 $pos=1 $flip=1
Mcpp incp incpb vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07 $pos=1 $flip=1
MI4 net52 incpb vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07 $pos=3 $flip=1
MI7 net85 incp vdd vdd sg13_lv_pmos l=1.300e-07 w=8.100e-07 $pos=3 $flip=1
Mdd0n d0 d net52 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07 $pos=4 $flip=1
Mdd0p d0 d net85 vdd sg13_lv_pmos l=1.300e-07 w=8.100e-07 $pos=4 $flip=1
MI47 d0 incp net59 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=5 $flip=0
MI45 d0 incpb net98 vdd sg13_lv_pmos l=1.300e-07 w=3.300e-07 $pos=5 $flip=0
MI48 net59 d1 net62 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=6 $flip=0
MI43 net98 d1 vdd vdd sg13_lv_pmos l=1.300e-07 w=3.050e-07 $pos=6 $flip=0
Mcdn0n net62 cdn vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=7 $flip=0
Md0d1n d1 d0 vss vss sg13_lv_nmos l=1.300e-07 w=4.300e-07 $pos=8 $flip=1
Mcdn0p net98 cdn vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07 $pos=8 $flip=0
Mswd1d2n d1 incp d2 vss sg13_lv_nmos l=1.300e-07 w=4.900e-07 $pos=9 $flip=0
Mdod1p d1 d0 vdd vdd sg13_lv_pmos l=1.300e-07 w=7.150e-07 $pos=9 $flip=1
MI23 d2 incpb net57 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=10 $flip=0
Mswd1d2p d1 incpb d2 vdd sg13_lv_pmos l=1.300e-07 w=1.030e-06 $pos=10 $flip=0
MI26 d2 incp net88 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07 $pos=11 $flip=0
MI24 net57 d3 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=12 $flip=0
MI28 net88 d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07 $pos=12 $flip=0
Mcdn1n net37 cdn vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07 $pos=13 $flip=1
Mcdn1p d3 cdn vdd vdd sg13_lv_pmos l=1.300e-07 w=9.900e-07 $pos=13 $flip=1
Md2d3n d3 d2 net37 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07 $pos=14 $flip=1
Md2d3p d3 d2 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.900e-07 $pos=14 $flip=0
Mobp q d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06 $pos=15 $flip=1
Mobn q d3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07 $pos=16 $flip=1
.ENDS


******* EOF

** Created by: circuit_gen.DFQD1_1
** Cell name: DFQD1_1
** Lib name: sg13g2
.SUBCKT sg13g2_DFQD1_1 cp d q vdd vss
*.PININFO cp:I d:I q:O vdd:B vss:B 
MI4 net43 incpb vss vss sg13_lv_nmos l=1.300e-07 w=4.050e-07
MI23 d2 incpb net42 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI5 d0 d net43 vss sg13_lv_nmos l=1.300e-07 w=4.050e-07
MI47 d0 incp net50 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI48 net50 d1 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI24 net42 d3 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI50 d1 incp d2 vss sg13_lv_nmos l=1.300e-07 w=3.750e-07
MI32_M_u2 incp incpb vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI31_M_u2 incpb cp vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI27_M_u2 q d3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI53_M_u2 d3 d2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI13_M_u2 d1 d0 vss vss sg13_lv_nmos l=1.300e-07 w=4.550e-07
MI6 d0 d net66 vdd sg13_lv_pmos l=1.300e-07 w=6.900e-07
MI32_M_u3 incp incpb vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI31_M_u3 incpb cp vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI27_M_u3 q d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI53_M_u3 d3 d2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI13_M_u3 d1 d0 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.900e-07
MI7 net66 incp vdd vdd sg13_lv_pmos l=1.300e-07 w=8.100e-07
MI52 d1 incpb d2 vdd sg13_lv_pmos l=1.300e-07 w=9.750e-07
MI28 net74 d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI26 d2 incp net74 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI45 d0 incpb net84 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI43 net84 d1 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
.ENDS


******* EOF

** Created by: circuit_gen.DFQD1_2
** Cell name: DFQD1_2
** Lib name: sg13g2
.SUBCKT sg13g2_DFQD1_2 cp d q vdd vss
*.PININFO cp:I d:I q:O vdd:B vss:B 
MI4 net43 incpb vss vss sg13_lv_nmos l=1.300e-07 w=4.050e-07
MI23 d2 incpb net42 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI5 d0 d net43 vss sg13_lv_nmos l=1.300e-07 w=4.050e-07
MI47 d0 incp net50 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI48 net50 d1 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI24 net42 d3 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI50 d1 incp d2 vss sg13_lv_nmos l=1.300e-07 w=3.750e-07
MI32_M_u2 incp incpb vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI31_M_u2 incpb cp vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI27_M_u2 q d3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI53_M_u2 d3 d2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI13_M_u2 d1 d0 vss vss sg13_lv_nmos l=1.300e-07 w=4.550e-07
MI6 d0 d net66 vdd sg13_lv_pmos l=1.300e-07 w=6.900e-07
MI32_M_u3 incp incpb vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI31_M_u3 incpb cp vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI27_M_u3 q d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI53_M_u3 d3 d2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI13_M_u3 d1 d0 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.900e-07
MI7 net66 incp vdd vdd sg13_lv_pmos l=1.300e-07 w=8.100e-07
MI52 d1 incpb d2 vdd sg13_lv_pmos l=1.300e-07 w=9.750e-07
MI28 net74 d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI26 d2 incp net74 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI45 d0 incpb net84 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI43 net84 d1 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
.ENDS


******* EOF

** Created by: circuit_gen.DFQD1_3
** Cell name: DFQD1_3
** Lib name: sg13g2
.SUBCKT sg13g2_DFQD1_3 cp d q vdd vss
*.PININFO cp:I d:I q:O vdd:B vss:B 
MI4 net43 incpb vss vss sg13_lv_nmos l=1.300e-07 w=4.050e-07
MI23 d2 incpb net42 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI5 d0 d net43 vss sg13_lv_nmos l=1.300e-07 w=4.050e-07
MI47 d0 incp net50 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI48 net50 d1 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI24 net42 d3 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI50 d1 incp d2 vss sg13_lv_nmos l=1.300e-07 w=3.750e-07
MI32_M_u2 incp incpb vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI31_M_u2 incpb cp vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI27_M_u2 q d3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI53_M_u2 d3 d2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI13_M_u2 d1 d0 vss vss sg13_lv_nmos l=1.300e-07 w=4.550e-07
MI6 d0 d net66 vdd sg13_lv_pmos l=1.300e-07 w=6.900e-07
MI32_M_u3 incp incpb vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI31_M_u3 incpb cp vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI27_M_u3 q d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI53_M_u3 d3 d2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI13_M_u3 d1 d0 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.900e-07
MI7 net66 incp vdd vdd sg13_lv_pmos l=1.300e-07 w=8.100e-07
MI52 d1 incpb d2 vdd sg13_lv_pmos l=1.300e-07 w=9.750e-07
MI28 net74 d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI26 d2 incp net74 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI45 d0 incpb net84 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI43 net84 d1 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
.ENDS


******* EOF

** Created by: circuit_gen.DFQD1
** Cell name: DFQD1
** Lib name: sg13g2
.SUBCKT sg13g2_DFQD1 cp d q vdd vss
*.PININFO cp:I d:I q:O vdd:B vss:B 
MI4 net43 incpb vss vss sg13_lv_nmos l=1.300e-07 w=4.050e-07
MI23 d2 incpb net42 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI5 d0 d net43 vss sg13_lv_nmos l=1.300e-07 w=4.050e-07
MI47 d0 incp net50 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI48 net50 d1 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI24 net42 d3 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
MI50 d1 incp d2 vss sg13_lv_nmos l=1.300e-07 w=3.750e-07
MI32_M_u2 incp incpb vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI31_M_u2 incpb cp vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI27_M_u2 q d3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI53_M_u2 d3 d2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI13_M_u2 d1 d0 vss vss sg13_lv_nmos l=1.300e-07 w=4.550e-07
MI6 d0 d net66 vdd sg13_lv_pmos l=1.300e-07 w=6.900e-07
MI32_M_u3 incp incpb vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI31_M_u3 incpb cp vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI27_M_u3 q d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI53_M_u3 d3 d2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI13_M_u3 d1 d0 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.900e-07
MI7 net66 incp vdd vdd sg13_lv_pmos l=1.300e-07 w=8.100e-07
MI52 d1 incpb d2 vdd sg13_lv_pmos l=1.300e-07 w=9.750e-07
MI28 net74 d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI26 d2 incp net74 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI45 d0 incpb net84 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
MI43 net84 d1 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07
.ENDS


******* EOF

** Created by: circuit_gen.FILL1
** Cell name: FILL1
** Lib name: sg13g2
.SUBCKT sg13g2_FILL1 vdd vss
*.PININFO vdd:B vss:B 
.ENDS


******* EOF

** Created by: circuit_gen.FILL2
** Cell name: FILL2
** Lib name: sg13g2
.SUBCKT sg13g2_FILL2 vdd vss
*.PININFO vdd:B vss:B 
.ENDS


******* EOF

** Created by: circuit_gen.FILL4
** Cell name: FILL4
** Lib name: sg13g2
.SUBCKT sg13g2_FILL4 vdd vss
*.PININFO vdd:B vss:B 
.ENDS


******* EOF

** Created by: circuit_gen.FILL8
** Cell name: FILL8
** Lib name: sg13g2
.SUBCKT sg13g2_FILL8 vdd vss
*.PININFO vdd:B vss:B 
.ENDS


******* EOF

** Created by: circuit_gen.INVD1_1
** Cell name: INVD1_1
** Lib name: sg13g2
.SUBCKT sg13g2_INVD1_1 i z vss vdd
*.PININFO i:I z:O vss:B vdd:B
M0 z i vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M1 z i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.INVD1_2
** Cell name: INVD1_2
** Lib name: sg13g2
.SUBCKT sg13g2_INVD1_2 i z vss vdd
*.PININFO i:I z:O vss:B vdd:B
M0 z i vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M1 z i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.INVD1_3
** Cell name: INVD1_3
** Lib name: sg13g2
.SUBCKT sg13g2_INVD1_3 i z vss vdd
*.PININFO i:I z:O vss:B vdd:B
M0 z i vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M1 z i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.INVD1
** Cell name: INVD1
** Lib name: sg13g2
.SUBCKT sg13g2_INVD1 i z vss vdd
*.PININFO i:I z:O vss:B vdd:B
M0 z i vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M1 z i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.MUX2D1_1
** Cell name: MUX2D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_MUX2D1_1 i0 i1 s vdd vss z
*.PININFO i0:I i1:I s:I z:O vdd:B vss:B 
MI15_M_u3 net46 s net28 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MU7_M_u3 net48 net42 net28 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI20_M_u2 net46 i1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI19_M_u2 net48 i0 vss vss sg13_lv_nmos l=1.300e-07 w=5.050e-07
MI18_M_u2 net42 s vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MU29_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI15_M_u2 net46 net42 net28 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MU7_M_u2 net48 s net28 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI20_M_u3 net46 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI19_M_u3 net48 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.100e-07
MI18_M_u3 net42 s vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MU29_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=7.700e-07
.ENDS


******* EOF

** Created by: circuit_gen.MUX2D1_2
** Cell name: MUX2D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_MUX2D1_2 i0 i1 s vdd vss z
*.PININFO i0:I i1:I s:I z:O vdd:B vss:B 
MI15_M_u3 net46 s net28 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MU7_M_u3 net48 net42 net28 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI20_M_u2 net46 i1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI19_M_u2 net48 i0 vss vss sg13_lv_nmos l=1.300e-07 w=5.050e-07
MI18_M_u2 net42 s vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MU29_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI15_M_u2 net46 net42 net28 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MU7_M_u2 net48 s net28 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI20_M_u3 net46 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI19_M_u3 net48 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.100e-07
MI18_M_u3 net42 s vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MU29_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=7.700e-07
.ENDS


******* EOF

** Created by: circuit_gen.MUX2D1_3
** Cell name: MUX2D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_MUX2D1_3 i0 i1 s vdd vss z
*.PININFO i0:I i1:I s:I z:O vdd:B vss:B 
MI15_M_u3 net46 s net28 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MU7_M_u3 net48 net42 net28 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI20_M_u2 net46 i1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI19_M_u2 net48 i0 vss vss sg13_lv_nmos l=1.300e-07 w=5.050e-07
MI18_M_u2 net42 s vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MU29_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI15_M_u2 net46 net42 net28 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MU7_M_u2 net48 s net28 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI20_M_u3 net46 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI19_M_u3 net48 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.100e-07
MI18_M_u3 net42 s vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MU29_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=7.700e-07
.ENDS


******* EOF

** Created by: circuit_gen.MUX2D1
** Cell name: MUX2D1
** Lib name: sg13g2
.SUBCKT sg13g2_MUX2D1 i0 i1 s vdd vss z
*.PININFO i0:I i1:I s:I z:O vdd:B vss:B 
MI15_M_u3 net46 s net28 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MU7_M_u3 net48 net42 net28 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI20_M_u2 net46 i1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI19_M_u2 net48 i0 vss vss sg13_lv_nmos l=1.300e-07 w=5.050e-07
MI18_M_u2 net42 s vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MU29_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI15_M_u2 net46 net42 net28 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MU7_M_u2 net48 s net28 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI20_M_u3 net46 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI19_M_u3 net48 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.100e-07
MI18_M_u3 net42 s vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MU29_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=7.700e-07
.ENDS


******* EOF

** Created by: circuit_gen.ND2D1_1
** Cell name: ND2D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_ND2D1_1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u3 zn a1 xi1_net6 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u4 xi1_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND2D1_2
** Cell name: ND2D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_ND2D1_2 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u3 zn a1 xi1_net6 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u4 xi1_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND2D1_3
** Cell name: ND2D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_ND2D1_3 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u3 zn a1 xi1_net6 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u4 xi1_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND2D1
** Cell name: ND2D1
** Lib name: sg13g2
.SUBCKT sg13g2_ND2D1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u3 zn a1 xi1_net6 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u4 xi1_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND3D1_1
** Cell name: ND3D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_ND3D1_1 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 xi1_net10 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u5 xi1_net10 a2 xi1_net13 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u6 xi1_net13 a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u3 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND3D1_2
** Cell name: ND3D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_ND3D1_2 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 xi1_net10 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u5 xi1_net10 a2 xi1_net13 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u6 xi1_net13 a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u3 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND3D1_3
** Cell name: ND3D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_ND3D1_3 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 xi1_net10 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u5 xi1_net10 a2 xi1_net13 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u6 xi1_net13 a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u3 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND3D1
** Cell name: ND3D1
** Lib name: sg13g2
.SUBCKT sg13g2_ND3D1 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 xi1_net10 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u5 xi1_net10 a2 xi1_net13 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u6 xi1_net13 a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u3 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND4D1_1
** Cell name: ND4D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_ND4D1_1 a1 a2 a3 a4 vdd vss zn
*.PININFO a1:I a2:I a3:I a4:I zn:O vdd:B vss:B 
MI3 p0 a2 p1 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI5 p2 a4 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4 p1 a3 p2 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MU53 zn a1 p0 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI7 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI2 zn a4 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI0 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND4D1_2
** Cell name: ND4D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_ND4D1_2 a1 a2 a3 a4 vdd vss zn
*.PININFO a1:I a2:I a3:I a4:I zn:O vdd:B vss:B 
MI3 p0 a2 p1 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI5 p2 a4 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4 p1 a3 p2 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MU53 zn a1 p0 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI7 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI2 zn a4 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI0 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND4D1_3
** Cell name: ND4D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_ND4D1_3 a1 a2 a3 a4 vdd vss zn
*.PININFO a1:I a2:I a3:I a4:I zn:O vdd:B vss:B 
MI3 p0 a2 p1 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI5 p2 a4 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4 p1 a3 p2 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MU53 zn a1 p0 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI7 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI2 zn a4 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI0 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.ND4D1
** Cell name: ND4D1
** Lib name: sg13g2
.SUBCKT sg13g2_ND4D1 a1 a2 a3 a4 vdd vss zn
*.PININFO a1:I a2:I a3:I a4:I zn:O vdd:B vss:B 
MI3 p0 a2 p1 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI5 p2 a4 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4 p1 a3 p2 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MU53 zn a1 p0 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI7 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI2 zn a4 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI0 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.NR2D1_1
** Cell name: NR2D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_NR2D1_1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u2 zn a1 xi1_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 xi1_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.NR2D1_2
** Cell name: NR2D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_NR2D1_2 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u2 zn a1 xi1_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 xi1_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.NR2D1_3
** Cell name: NR2D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_NR2D1_3 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u2 zn a1 xi1_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 xi1_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.NR2D1
** Cell name: NR2D1
** Lib name: sg13g2
.SUBCKT sg13g2_NR2D1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI1_M_u2 zn a1 xi1_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI1_M_u1 xi1_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.NR3D1_1
** Cell name: NR3D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_NR3D1_1 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
M_u4 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI2 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI3 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4_0 net37_0_ a2 net34_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u1_0 net34_0_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u1_1 net34_1_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI4_1 net37_1_ a2 net34_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_0 zn a1 net37_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_1 zn a1 net37_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.NR3D1_2
** Cell name: NR3D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_NR3D1_2 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
M_u4 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI2 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI3 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4_0 net37_0_ a2 net34_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u1_0 net34_0_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u1_1 net34_1_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI4_1 net37_1_ a2 net34_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_0 zn a1 net37_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_1 zn a1 net37_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.NR3D1_3
** Cell name: NR3D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_NR3D1_3 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
M_u4 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI2 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI3 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4_0 net37_0_ a2 net34_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u1_0 net34_0_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u1_1 net34_1_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI4_1 net37_1_ a2 net34_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_0 zn a1 net37_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_1 zn a1 net37_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.NR3D1
** Cell name: NR3D1
** Lib name: sg13g2
.SUBCKT sg13g2_NR3D1 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
M_u4 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI2 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI3 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4_0 net37_0_ a2 net34_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u1_0 net34_0_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u1_1 net34_1_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI4_1 net37_1_ a2 net34_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_0 zn a1 net37_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_1 zn a1 net37_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OA21D1_1
** Cell name: OA21D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_OA21D1_1 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI12 net14 a2 net20 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI11 net14 a1 net20 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI6 net20 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI8_M_u2 z net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI9 net14 a1 net24 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI8_M_u3 z net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net14 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI7 net24 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OA21D1_2
** Cell name: OA21D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_OA21D1_2 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI12 net14 a2 net20 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI11 net14 a1 net20 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI6 net20 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI8_M_u2 z net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI9 net14 a1 net24 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI8_M_u3 z net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net14 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI7 net24 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OA21D1_3
** Cell name: OA21D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_OA21D1_3 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI12 net14 a2 net20 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI11 net14 a1 net20 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI6 net20 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI8_M_u2 z net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI9 net14 a1 net24 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI8_M_u3 z net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net14 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI7 net24 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OA21D1
** Cell name: OA21D1
** Lib name: sg13g2
.SUBCKT sg13g2_OA21D1 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI12 net14 a2 net20 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI11 net14 a1 net20 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI6 net20 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI8_M_u2 z net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI9 net14 a1 net24 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI8_M_u3 z net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u2 net14 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI7 net24 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OAI21D1_1
** Cell name: OAI21D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_OAI21D1_1 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
M_u2 zn a1 net15 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u3 zn a2 net15 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u4 net15 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI16_MI12 zn a1 xi16_net11 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u9 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI16_MI13 xi16_net11 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OAI21D1_2
** Cell name: OAI21D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_OAI21D1_2 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
M_u2 zn a1 net15 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u3 zn a2 net15 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u4 net15 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI16_MI12 zn a1 xi16_net11 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u9 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI16_MI13 xi16_net11 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OAI21D1_3
** Cell name: OAI21D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_OAI21D1_3 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
M_u2 zn a1 net15 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u3 zn a2 net15 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u4 net15 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI16_MI12 zn a1 xi16_net11 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u9 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI16_MI13 xi16_net11 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OAI21D1
** Cell name: OAI21D1
** Lib name: sg13g2
.SUBCKT sg13g2_OAI21D1 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
M_u2 zn a1 net15 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u3 zn a2 net15 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u4 net15 b vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI16_MI12 zn a1 xi16_net11 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u9 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI16_MI13 xi16_net11 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OR2D1_1
** Cell name: OR2D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_OR2D1_1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MU1_M_u2 z net7 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u4 net7 a1 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u3 net7 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u2 net7 a1 x_u7_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MU1_M_u3 z net7 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u7_M_u1 x_u7_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OR2D1_2
** Cell name: OR2D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_OR2D1_2 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MU1_M_u2 z net7 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u4 net7 a1 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u3 net7 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u2 net7 a1 x_u7_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MU1_M_u3 z net7 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u7_M_u1 x_u7_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OR2D1_3
** Cell name: OR2D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_OR2D1_3 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MU1_M_u2 z net7 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u4 net7 a1 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u3 net7 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u2 net7 a1 x_u7_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MU1_M_u3 z net7 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u7_M_u1 x_u7_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.OR2D1
** Cell name: OR2D1
** Lib name: sg13g2
.SUBCKT sg13g2_OR2D1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MU1_M_u2 z net7 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u4 net7 a1 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u3 net7 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.350e-07
M_u7_M_u2 net7 a1 x_u7_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MU1_M_u3 z net7 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u7_M_u1 x_u7_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.TAPCELL
** Cell name: TAPCELL
** Lib name: sg13g2
.SUBCKT sg13g2_TAPCELL vdd vss
*.PININFO vdd:B vss:B 
.ENDS


******* EOF

** Created by: circuit_gen.TIEH_1
** Cell name: TIEH_1
** Lib name: sg13g2
.SUBCKT sg13g2_TIEH_1 vdd vss z
*.PININFO z:O vdd:B vss:B 
M_u2 net6 net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u1 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.TIEH_2
** Cell name: TIEH_2
** Lib name: sg13g2
.SUBCKT sg13g2_TIEH_2 vdd vss z
*.PININFO z:O vdd:B vss:B 
M_u2 net6 net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u1 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.TIEH_3
** Cell name: TIEH_3
** Lib name: sg13g2
.SUBCKT sg13g2_TIEH_3 vdd vss z
*.PININFO z:O vdd:B vss:B 
M_u2 net6 net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u1 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.TIEH
** Cell name: TIEH
** Lib name: sg13g2
.SUBCKT sg13g2_TIEH vdd vss z
*.PININFO z:O vdd:B vss:B 
M_u2 net6 net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u1 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.TIEL_1
** Cell name: TIEL_1
** Lib name: sg13g2
.SUBCKT sg13g2_TIEL_1 vdd vss zn
*.PININFO zn:O vdd:B vss:B 
M_u2 zn net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u1 net6 net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.TIEL_2
** Cell name: TIEL_2
** Lib name: sg13g2
.SUBCKT sg13g2_TIEL_2 vdd vss zn
*.PININFO zn:O vdd:B vss:B 
M_u2 zn net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u1 net6 net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.TIEL_3
** Cell name: TIEL_3
** Lib name: sg13g2
.SUBCKT sg13g2_TIEL_3 vdd vss zn
*.PININFO zn:O vdd:B vss:B 
M_u2 zn net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u1 net6 net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.TIEL
** Cell name: TIEL
** Lib name: sg13g2
.SUBCKT sg13g2_TIEL vdd vss zn
*.PININFO zn:O vdd:B vss:B 
M_u2 zn net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u1 net6 net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
.ENDS


******* EOF

** Created by: circuit_gen.XNR2D1_1
** Cell name: XNR2D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_XNR2D1_1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
M_u2_M_u2 net4 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u5_M_u2 net6 net4 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u4_M_u2 zn net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u8_M_u2 net10 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u6_M_u3 net4 a1 net14 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u7_M_u3 net6 net10 net14 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u6_M_u2 net4 net10 net14 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u2_M_u3 net4 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u5_M_u3 net6 net4 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u4_M_u3 zn net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u8_M_u3 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u7_M_u2 net6 a1 net14 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.XNR2D1_2
** Cell name: XNR2D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_XNR2D1_2 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
M_u2_M_u2 net4 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u5_M_u2 net6 net4 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u4_M_u2 zn net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u8_M_u2 net10 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u6_M_u3 net4 a1 net14 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u7_M_u3 net6 net10 net14 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u6_M_u2 net4 net10 net14 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u2_M_u3 net4 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u5_M_u3 net6 net4 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u4_M_u3 zn net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u8_M_u3 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u7_M_u2 net6 a1 net14 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.XNR2D1_3
** Cell name: XNR2D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_XNR2D1_3 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
M_u2_M_u2 net4 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u5_M_u2 net6 net4 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u4_M_u2 zn net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u8_M_u2 net10 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u6_M_u3 net4 a1 net14 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u7_M_u3 net6 net10 net14 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u6_M_u2 net4 net10 net14 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u2_M_u3 net4 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u5_M_u3 net6 net4 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u4_M_u3 zn net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u8_M_u3 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u7_M_u2 net6 a1 net14 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.XNR2D1
** Cell name: XNR2D1
** Lib name: sg13g2
.SUBCKT sg13g2_XNR2D1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
M_u2_M_u2 net4 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u5_M_u2 net6 net4 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u4_M_u2 zn net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
M_u8_M_u2 net10 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u6_M_u3 net4 a1 net14 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u7_M_u3 net6 net10 net14 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
M_u6_M_u2 net4 net10 net14 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u2_M_u3 net4 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u5_M_u3 net6 net4 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u4_M_u3 zn net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
M_u8_M_u3 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
M_u7_M_u2 net6 a1 net14 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.XOR2D1_1
** Cell name: XOR2D1_1
** Lib name: sg13g2
.SUBCKT sg13g2_XOR2D1_1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MI6_M_u3 net41 a1 net21 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI2_M_u3 net27 net23 net21 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI7_M_u2 net41 net27 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI3_M_u2 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4_M_u2 z net21 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI5_M_u2 net23 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI6_M_u2 net41 net23 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI2_M_u2 net27 a1 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI7_M_u3 net41 net27 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI3_M_u3 net27 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI4_M_u3 z net21 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_M_u3 net23 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.XOR2D1_2
** Cell name: XOR2D1_2
** Lib name: sg13g2
.SUBCKT sg13g2_XOR2D1_2 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MI6_M_u3 net41 a1 net21 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI2_M_u3 net27 net23 net21 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI7_M_u2 net41 net27 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI3_M_u2 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4_M_u2 z net21 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI5_M_u2 net23 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI6_M_u2 net41 net23 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI2_M_u2 net27 a1 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI7_M_u3 net41 net27 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI3_M_u3 net27 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI4_M_u3 z net21 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_M_u3 net23 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.XOR2D1_3
** Cell name: XOR2D1_3
** Lib name: sg13g2
.SUBCKT sg13g2_XOR2D1_3 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MI6_M_u3 net41 a1 net21 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI2_M_u3 net27 net23 net21 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI7_M_u2 net41 net27 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI3_M_u2 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4_M_u2 z net21 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI5_M_u2 net23 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI6_M_u2 net41 net23 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI2_M_u2 net27 a1 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI7_M_u3 net41 net27 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI3_M_u3 net27 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI4_M_u3 z net21 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_M_u3 net23 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

** Created by: circuit_gen.XOR2D1
** Cell name: XOR2D1
** Lib name: sg13g2
.SUBCKT sg13g2_XOR2D1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MI6_M_u3 net41 a1 net21 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI2_M_u3 net27 net23 net21 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI7_M_u2 net41 net27 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI3_M_u2 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI4_M_u2 z net21 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07
MI5_M_u2 net23 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07
MI6_M_u2 net41 net23 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI2_M_u2 net27 a1 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI7_M_u3 net41 net27 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
MI3_M_u3 net27 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI4_M_u3 z net21 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06
MI5_M_u3 net23 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07
.ENDS


******* EOF

************************************************************************
* Customized version of the sg13g2_io because the LVS is trash
* Put the sub pin in order to be connected to VSS later, as god intended
* It would be helpful if there is a way to check LVS with IO and pads 
* without so much trouble
************************************************************************

************************************************************************
*
* Copyright 2024 IHP PDK Authors
* 
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
* 
*    https://www.apache.org/licenses/LICENSE-2.0
* 
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

**ptap1 (TIE SUB)
.subckt ptap1 1 2 r=22.472 A=24.01p Perim=19.6u w=4.9u l=4.9u
* TODO: The LVS (up to aug/28) doesnt extract correctly
*       or extracts correctly, but cannot merge/compare
*R1 1 2 R=r A=A P=Perim w=w l=l
*D1 2 1 ptap1 A=A P=Perim
.ends ptap1

**ntap1 (TIE WELL)
.subckt ntap1 1 2 r=22.472 A=24.01p Perim=19.6u w=4.9u l=4.9u
* TODO: The LVS (up to aug/28) doesnt extract correctly
*       or extracts correctly, but cannot merge/compare
*R1 1 2 R=r A=A P=Perim w=w l=l
*D1 1 2 ntap1 A=A P=Perim
.ends ntap1

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadIOVss
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadIOVss iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
DD4 sub iovss dantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
DD2 sub iovss dantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
DD3 iovss iovdd dpantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
DD1 iovss iovdd dpantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
XR2 vss sub / ptap1 r=22.472 A=24.01p Perim=19.6u w=4.9u l=4.9u
XR0 iovss sub / ptap1 r=169.45m A=5.487n Perim=296.3u w=74.075u l=74.075u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_N43N43D4R
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_N43N43D4R gate pad tie sub
*.PININFO gate:I pad:B tie:B
MN0<1> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<2> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<3> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<4> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<5> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<6> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<7> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<8> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<9> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<10> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<11> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<12> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<13> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<14> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<15> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<16> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<17> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<18> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<19> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<20> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<21> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<22> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<23> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<24> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<25> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<26> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<27> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<28> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<29> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<30> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<31> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<32> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<33> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<34> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<35> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<36> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<37> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<38> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<39> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<40> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<41> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<42> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<43> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<44> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<45> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<46> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<47> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<48> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<49> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<50> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<51> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<52> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<53> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<54> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<55> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<56> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<57> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<58> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<59> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<60> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<61> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<62> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<63> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<64> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<65> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<66> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<67> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<68> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<69> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<70> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<71> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<72> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<73> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<74> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<75> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<76> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<77> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<78> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<79> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<80> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<81> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<82> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<83> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<84> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<85> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<86> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<87> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<88> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<89> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<90> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<91> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<92> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<93> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<94> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<95> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<96> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<97> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<98> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<99> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<100> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<101> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<102> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<103> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<104> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<105> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<106> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<107> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<108> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<109> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<110> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<111> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<112> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<113> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<114> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<115> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<116> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<117> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<118> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<119> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<120> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<121> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<122> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<123> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<124> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<125> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<126> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<127> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<128> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<129> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<130> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<131> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<132> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<133> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<134> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<135> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<136> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<137> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<138> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<139> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<140> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<141> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<142> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<143> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<144> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<145> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<146> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<147> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<148> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<149> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<150> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<151> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<152> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<153> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<154> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<155> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<156> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<157> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<158> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<159> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<160> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<161> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<162> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<163> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<164> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<165> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<166> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<167> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<168> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<169> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<170> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<171> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<172> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
XR0 tie sub / ptap1 r=9.999 A=65.61p Perim=32.4u w=8.1u l=8.1u
DD0 sub gate dantenna m=1 w=480n l=480n a=230.4f p=1.92u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_RCClampResistor
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_RCClampResistor pin1 pin2 sub
*.PININFO pin1:B pin2:B
R$274 pin2 pin1 rppd w=1u l=520u ps=0 b=0 m=1
*RR29 net15 net16 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR28 net20 net21 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR27 net23 net24 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR24 net17 net18 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR23 net16 net17 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR21 net25 pin2 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR20 net22 net23 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR19 net19 net20 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR17 net24 net25 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR16 net21 net22 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR15 net18 net19 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR14 net5 net6 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR13 net8 net9 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR12 net11 net12 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR11 net14 net15 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR10 net2 net3 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR9 net1 net2 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
*RR8 net13 net14 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR7 net10 net11 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR6 net7 net8 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
*RR5 net4 net5 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
*RR4 net12 net13 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR3 net9 net10 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
*+ b=0
*RR2 net6 net7 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
*RR1 net3 net4 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
*RR0 pin1 net1 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_RCClampInverter
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_RCClampInverter in iovss out supply sub
*.PININFO in:B iovss:B out:B supply:B
MN1 iovss in iovss sub sg13_hv_nmos m=1 w=126.000u l=9.5u ng=14
MN0 out in iovss sub sg13_hv_nmos m=1 w=108.000u l=500.0n ng=12
XR0 iovss sub / ptap1 r=9.59 A=68.973p Perim=33.22u w=8.305u l=8.305u
MP0 out in supply supply sg13_hv_pmos m=1 w=350.000u l=500.0n ng=50
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadVdd
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadVdd iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XI0 net2 vdd iovss sub / sg13g2_Clamp_N43N43D4R
XI2 vdd net1 sub / sg13g2_RCClampResistor
XR1 iovss sub / ptap1 r=456.33m A=1.97n Perim=177.54u w=44.385u l=44.385u
XR0 vss sub / ptap1 r=22.472 A=24.01p Perim=19.6u w=4.9u l=4.9u
XI1 net1 iovss net2 vdd sub / sg13g2_RCClampInverter
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadIOVdd
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadIOVdd iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XI0 net2 iovdd iovss sub / sg13g2_Clamp_N43N43D4R
XI2 iovdd net1 sub / sg13g2_RCClampResistor
XI1 net1 iovss net2 iovdd sub / sg13g2_RCClampInverter
XR1 iovss sub / ptap1 r=449.797m A=2n Perim=178.88u w=44.72u l=44.72u
XR0 vss sub / ptap1 r=22.832 A=23.523p Perim=19.4u w=4.85u l=4.85u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_DCNDiode
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_DCNDiode anode cathode guard sub
*.PININFO anode:B cathode:B guard:B
DD1 sub cathode dantenna m=1 w=1.26u l=27.78u a=35.0028p p=58.08u
DD0 sub cathode dantenna m=1 w=1.26u l=27.78u a=35.0028p p=58.08u
*XR0 anode sub / ptap1 r=5.191 A=141.253p Perim=47.54u w=11.885u l=11.885u
XR0 anode sub / ptap1 r=5.191 A=141.2964p Perim=221.76u w=11.885u l=11.885u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_DCPDiode
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_DCPDiode anode cathode guard sub
*.PININFO anode:B cathode:B guard:B
DD1 anode cathode dpantenna m=1 w=1.26u l=27.78u a=35.0028p p=58.08u
DD0 anode cathode dpantenna m=1 w=1.26u l=27.78u a=35.0028p p=58.08u
*XR0 guard sub / ptap1 r=17.289 A=33.524p Perim=23.16u w=5.79u l=5.79u
XR0 guard sub / ptap1 r=17.289 A=33.5104p Perim=197.12u w=5.79u l=5.79u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadVss
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadVss iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XI1 iovss vss iovss sub / sg13g2_DCNDiode
XI2 vss iovdd iovss sub / sg13g2_DCPDiode
XR1 iovss sub / ptap1 r=174.346m A=5.329n Perim=292u w=73u l=73u
XR0 vss sub / ptap1 r=22.832 A=23.523p Perim=19.4u w=4.85u l=4.85u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Filler4000
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Filler4000 iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XR1 vss sub / ptap1 r=63.078 A=5.856p Perim=9.68u w=2.42u l=2.42u
XR0 iovss sub / ptap1 r=625.742m A=1.416n Perim=150.5u w=37.625u l=37.625u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_io_inv_x1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_io_inv_x1 i nq vdd vss sub
*.PININFO i:I nq:O vdd:B vss:B
MN0 nq i vss sub sg13_lv_nmos m=1 w=3.93u l=130.00n ng=1
MP0 nq i vdd vdd sg13_lv_pmos m=1 w=4.41u l=130.00n ng=1
XR0 vss sub / ptap1 r=258.978 A=624.1f Perim=3.16u w=790n l=790n
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_LevelUp
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_LevelUp i iovdd o vdd vss sub
*.PININFO i:I o:O iovdd:B vdd:B vss:B
MN0 net2 i vss sub sg13_lv_nmos m=1 w=2.75u l=130.00n ng=1
MP0 net2 i vdd vdd sg13_lv_pmos m=1 w=4.75u l=130.00n ng=1
MN3 o net4 vss sub sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MN2 net4 i vss sub sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MN1 net3 net2 vss sub sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MP3 o net4 iovdd iovdd sg13_hv_pmos m=1 w=3.9u l=450.00n ng=1
MP2 net3 net4 iovdd iovdd sg13_hv_pmos m=1 w=300.0n l=450.00n ng=1
MP1 net4 net3 iovdd iovdd sg13_hv_pmos m=1 w=300.0n l=450.00n ng=1
XR0 vss sub / ptap1 r=207.099 A=912.025f Perim=3.82u w=955n l=955n
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_io_nor2_x1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_io_nor2_x1 i0 i1 nq vdd vss sub
*.PININFO i0:I i1:I nq:O vdd:B vss:B
MN0 nq i0 vss sub sg13_lv_nmos m=1 w=3.93u l=130.00n ng=1
MN1 nq i1 vss sub sg13_lv_nmos m=1 w=3.93u l=130.00n ng=1
MP1 net1 i0 vdd vdd sg13_lv_pmos m=1 w=4.41u l=130.00n ng=1
MP0 nq i1 net1 vdd sg13_lv_pmos m=1 w=4.41u l=130.00n ng=1
XR0 vss sub / ptap1 r=251.534 A=656.1f Perim=3.24u w=810n l=810n
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_io_tie
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_io_tie vdd vss sub
*.PININFO vdd:B vss:B
XR0 vss sub / ptap1 r=258.978 A=624.1f Perim=3.16u w=790n l=790n
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_io_nand2_x1
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_io_nand2_x1 i0 i1 nq vdd vss sub
*.PININFO i0:I i1:I nq:O vdd:B vss:B
MP1 nq i1 vdd vdd sg13_lv_pmos m=1 w=4.41u l=130.00n ng=1
MP0 nq i0 vdd vdd sg13_lv_pmos m=1 w=4.41u l=130.00n ng=1
MN1 net1 i0 vss sub sg13_lv_nmos m=1 w=3.93u l=130.00n ng=1
MN0 nq i1 net1 sub sg13_lv_nmos m=1 w=3.93u l=130.00n ng=1
XR0 vss sub / ptap1 r=251.534 A=656.1f Perim=3.24u w=810n l=810n
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_GateDecode
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_GateDecode core en iovdd ngate pgate vdd vss sub
*.PININFO core:I en:I ngate:O pgate:O iovdd:B vdd:B vss:B
XI2 en net3 vdd vss sub / sg13g2_io_inv_x1
XI4 net4 iovdd ngate vdd vss sub / sg13g2_LevelUp
XI3 net2 iovdd pgate vdd vss sub / sg13g2_LevelUp
XI0 core net3 net4 vdd vss sub / sg13g2_io_nor2_x1
XI5 vdd vss sub / sg13g2_io_tie
XI1 core en net2 vdd vss sub / sg13g2_io_nand2_x1
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_N2N2D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_N2N2D gate iovss pad sub
*.PININFO gate:B iovss:B pad:B
XR0 iovss sub / ptap1 r=11.438 A=55.801p Perim=29.88u w=7.47u l=7.47u
MN1 iovss gate pad sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0 pad gate iovss sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
DD0 sub gate dantenna m=1 w=780.00n l=780.00n a=608.400f p=3.12u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_P2N2D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_P2N2D gate iovdd iovss pad sub
*.PININFO gate:B iovdd:B iovss:B pad:B
DD0 gate iovdd dpantenna m=1 w=480n l=480n a=230.4f p=1.92u
MP1 iovdd gate pad iovdd sg13_hv_pmos m=1 w=13.32u l=600.0n ng=2
MP0 pad gate iovdd iovdd sg13_hv_pmos m=1 w=13.32u l=600.0n ng=2
XR0 iovss sub / ptap1 r=9.826 A=66.994p Perim=32.74u w=8.185u l=8.185u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_SecondaryProtection
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_SecondaryProtection core minus pad plus sub
*.PININFO core:B minus:B pad:B plus:B
*RR0 pad core 586.899 $SUB=sub $[res_rppd] m=1 l=2u w=1u ps=180n trise=0.0 b=0
RR0 pad core rppd m=1 l=2u w=1u
DD0 sub core dantenna m=1 w=640n l=3.1u a=1.984p p=7.48u
*XR1 minus sub / ptap1 r=46.556 A=9.03p Perim=12.02u w=3.005u l=3.005u
XR1 minus sub / ptap1 r=46.556 A=9.0304p Perim=53.12u w=3.005u l=3.005u
DD1 core plus dpantenna m=1 w=640n l=4.98u a=3.187p p=11.24u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_LevelDown
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_LevelDown core iovdd iovss pad vdd vss sub
*.PININFO core:O iovdd:B iovss:B pad:B vdd:B vss:B
MP0 net2 net4 vdd vdd sg13_hv_pmos m=1 w=4.65u l=450.00n ng=1
MN0 net2 net4 vss sub sg13_hv_nmos m=1 w=2.65u l=450.00n ng=1
MN1 core net2 vss sub sg13_lv_nmos m=1 w=2.75u l=130.00n ng=1
MP1 core net2 vdd vdd sg13_lv_pmos m=1 w=4.75u l=130.00n ng=1
*XR0 vss sub / ptap1 r=127.332 A=2.016p Perim=5.68u w=1.42u l=1.42u
XR0 vss sub / ptap1 r=127.332 A=2.019p Perim=14.06u w=1.42u l=1.42u
XI0 net4 iovss pad iovdd sub / sg13g2_SecondaryProtection
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadInOut4mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadInOut4mA c2p c2p_en iovdd iovss p2c pad vdd vss sub
*.PININFO c2p:I c2p_en:I p2c:O iovdd:B iovss:B pad:B vdd:B vss:B
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XI0 c2p c2p_en iovdd net2 net1 vdd vss sub / sg13g2_GateDecode
XI7 net2 iovss pad sub / sg13g2_Clamp_N2N2D
XI6 net1 iovdd iovss pad sub / sg13g2_Clamp_P2N2D
XI1 p2c iovdd iovss pad vdd vss sub / sg13g2_LevelDown
XR1 vss sub / ptap1 r=26.933 A=18.966p Perim=17.42u w=4.355u l=4.355u
XR0 iovss sub / ptap1 r=214.134m A=4.314n Perim=262.72u w=65.68u l=65.68u
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_P15N15D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_P15N15D gate iovdd iovss pad sub
*.PININFO gate:B iovdd:B iovss:B pad:B
DD0 gate iovdd dpantenna m=1 w=780.00n l=780.00n a=608.400f p=3.12u
XR0 iovss sub / ptap1 r=9.826 A=66.994p Perim=32.74u w=8.185u l=8.185u
MP1 pad gate iovdd iovdd sg13_hv_pmos m=1 w=199.8u l=600.0n ng=30
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_N15N15D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_N15N15D gate iovss pad sub
*.PININFO gate:B iovss:B pad:B
XR0 iovss sub / ptap1 r=11.438 A=55.801p Perim=29.88u w=7.47u l=7.47u
MN0 pad gate iovss sub sg13_hv_nmos m=1 w=66.000u l=600.0n ng=15
DD0 sub gate dantenna m=1 w=780.00n l=780.00n a=608.400f p=3.12u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadInOut30mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadInOut30mA c2p c2p_en iovdd iovss p2c pad vdd vss sub
*.PININFO c2p:I c2p_en:I p2c:O iovdd:B iovss:B pad:B vdd:B vss:B
XI1 p2c iovdd iovss pad vdd vss sub / sg13g2_LevelDown
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XI7 net1 iovdd iovss pad sub / sg13g2_Clamp_P15N15D
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI6 net2 iovss pad sub / sg13g2_Clamp_N15N15D
XR4 vss sub / ptap1 r=26.746 A=19.141p Perim=17.5u w=4.375u l=4.375u
XR3 iovss sub / ptap1 r=214.165m A=4.313n Perim=262.7u w=65.675u l=65.675u
XI0 c2p c2p_en iovdd net2 net1 vdd vss sub / sg13g2_GateDecode
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_LevelUpInv
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_LevelUpInv i iovdd o vdd vss sub
*.PININFO i:I o:O iovdd:B vdd:B vss:B
MN0 net2 i vss sub sg13_lv_nmos m=1 w=2.75u l=130.00n ng=1
MP0 net2 i vdd vdd sg13_lv_pmos m=1 w=4.75u l=130.00n ng=1
MN3 o net4 vss sub sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MN2 net4 net2 vss sub sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MN1 net3 i vss sub sg13_hv_nmos m=1 w=1.9u l=450.00n ng=1
MP3 o net4 iovdd iovdd sg13_hv_pmos m=1 w=3.9u l=450.00n ng=1
MP2 net3 net4 iovdd iovdd sg13_hv_pmos m=1 w=300.0n l=450.00n ng=1
MP1 net4 net3 iovdd iovdd sg13_hv_pmos m=1 w=300.0n l=450.00n ng=1
XR0 vss sub / ptap1 r=190.268 A=1.051p Perim=4.1u w=1.025u l=1.025u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_GateLevelUpInv
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_GateLevelUpInv core iovdd ngate pgate vdd vss sub
*.PININFO core:I ngate:O pgate:O iovdd:B vdd:B vss:B
XI1 core iovdd pgate vdd vss sub / sg13g2_LevelUpInv
XI0 core iovdd ngate vdd vss sub / sg13g2_LevelUpInv
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadOut4mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadOut4mA c2p iovdd iovss pad vdd vss sub
*.PININFO c2p:I iovdd:B iovss:B pad:B vdd:B vss:B
XI6 c2p iovdd net2 net1 vdd vss sub / sg13g2_GateLevelUpInv
XI7 net1 iovdd iovss pad sub / sg13g2_Clamp_P2N2D
XI8 net2 iovss pad sub / sg13g2_Clamp_N2N2D
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XR2 iovss sub / ptap1 r=212.747m A=4.343n Perim=263.6u w=65.9u l=65.9u
XR1 vss sub / ptap1 r=24.125 A=21.902p Perim=18.72u w=4.68u l=4.68u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadOut30mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadOut30mA c2p iovdd iovss pad vdd vss sub
*.PININFO c2p:I iovdd:B iovss:B pad:B vdd:B vss:B
XI6 c2p iovdd net2 net1 vdd vss sub / sg13g2_GateLevelUpInv
XI7 net1 iovdd iovss pad sub / sg13g2_Clamp_P15N15D
XI8 net2 iovss pad sub / sg13g2_Clamp_N15N15D
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XR1 vss sub / ptap1 r=24.125 A=21.902p Perim=18.72u w=4.68u l=4.68u
XR2 iovss sub / ptap1 r=214.165m A=4.313n Perim=262.7u w=65.675u l=65.675u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadIn
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadIn iovdd iovss p2c pad vdd vss sub
.PININFO p2c:O iovdd:B iovss:B pad:B vdd:B vss:B
XI1 p2c iovdd iovss pad vdd vss sub / sg13g2_LevelDown
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
*XR1 vss sub / ptap1 r=24.69 A=21.252p Perim=18.44u w=4.61u l=4.61u
*XR2 iovss sub / ptap1 r=173.674m A=5.35n Perim=292.58u w=73.145u l=73.145u
XR1 vss sub / ptap1 r=24.69 A=21.981p Perim=107.48u w=4.61u l=4.61u
XR2 iovss sub / ptap1 r=173.674m A=5223.2628p Perim=221.16u w=73.145u l=73.145u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_P8N8D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_P8N8D gate iovdd iovss pad sub
*.PININFO gate:B iovdd:B iovss:B pad:B
XR0 iovss sub / ptap1 r=9.826 A=66.994p Perim=32.74u w=8.185u l=8.185u
MP0 pad gate iovdd iovdd sg13_hv_pmos m=1 w=106.56u l=600.0n ng=16
DD0 gate iovdd dpantenna m=1 w=480n l=480n a=230.4f p=1.92u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_N8N8D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_N8N8D gate iovss pad sub
*.PININFO gate:B iovss:B pad:B
XR0 iovss sub / ptap1 r=11.438 A=55.801p Perim=29.88u w=7.47u l=7.47u
MN0 pad gate iovss sub sg13_hv_nmos m=1 w=35.2u l=600.0n ng=8
DD0 sub gate dantenna m=1 w=780.00n l=780.00n a=608.400f p=3.12u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadInOut16mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadInOut16mA c2p c2p_en iovdd iovss p2c pad vdd vss sub
*.PININFO c2p:I c2p_en:I p2c:O iovdd:B iovss:B pad:B vdd:B vss:B
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XI0 c2p c2p_en iovdd net2 net1 vdd vss sub / sg13g2_GateDecode
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI7 net1 iovdd iovss pad sub / sg13g2_Clamp_P8N8D
XI1 p2c iovdd iovss pad vdd vss sub / sg13g2_LevelDown
XI6 net2 iovss pad sub / sg13g2_Clamp_N8N8D
XR1 vss sub / ptap1 r=26.933 A=18.966p Perim=17.42u w=4.355u l=4.355u
XR0 iovss sub / ptap1 r=207.756m A=4.45n Perim=266.84u w=66.71u l=66.71u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadOut16mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadOut16mA c2p iovdd iovss pad vdd vss sub
*.PININFO c2p:I iovdd:B iovss:B pad:B vdd:B vss:B
* TODO: AGAIN?!?!?!
*XI6 c2p iovdda net2 net1 vdd vss sub / sg13g2_GateLevelUpInv
XI6 c2p iovdd net2 net1 vdd vss sub / sg13g2_GateLevelUpInv
XI8 net1 iovdd iovss pad sub / sg13g2_Clamp_P8N8D
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI7 net2 iovss pad sub / sg13g2_Clamp_N8N8D
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XR1 vss sub / ptap1 r=23.888 A=22.184p Perim=18.84u w=4.71u l=4.71u
XR2 iovss sub / ptap1 r=208.667m A=4.43n Perim=266.24u w=66.56u l=66.56u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadTriOut4mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadTriOut4mA c2p c2p_en iovdd iovss pad vdd vss sub
*.PININFO c2p:I c2p_en:I iovdd:B iovss:B pad:B vdd:B vss:B
XI7 c2p c2p_en iovdd net2 net1 vdd vss sub / sg13g2_GateDecode
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI8 net2 iovss pad sub / sg13g2_Clamp_N2N2D
XI9 net1 iovdd iovss pad sub / sg13g2_Clamp_P2N2D
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XR1 vss sub / ptap1 r=24.567 A=21.391p Perim=18.5u w=4.625u l=4.625u
XR2 iovss sub / ptap1 r=208.667m A=4.43n Perim=266.24u w=66.56u l=66.56u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadTriOut16mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadTriOut16mA c2p c2p_en iovdd iovss pad vdd vss sub
*.PININFO c2p:I c2p_en:I iovdd:B iovss:B pad:B vdd:B vss:B
XI7 c2p c2p_en iovdd net2 net1 vdd vss sub / sg13g2_GateDecode
XI8 net1 iovdd iovss pad sub / sg13g2_Clamp_P8N8D
XI9 net2 iovss pad sub / sg13g2_Clamp_N8N8D
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XR1 vss sub / ptap1 r=24.897 A=21.022p Perim=18.34u w=4.585u l=4.585u
XR2 iovss sub / ptap1 r=208.211m A=4.44n Perim=266.54u w=66.635u l=66.635u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadTriOut30mA
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadTriOut30mA c2p c2p_en iovdd iovss pad vdd vss sub
*.PININFO c2p:I c2p_en:I iovdd:B iovss:B pad:B vdd:B vss:B
XI7 c2p c2p_en iovdd net2 net1 vdd vss sub / sg13g2_GateDecode
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI8 net2 iovss pad sub / sg13g2_Clamp_N15N15D
XI9 net1 iovdd iovss pad sub / sg13g2_Clamp_P15N15D
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
XR1 vss sub / ptap1 r=24.649 A=21.298p Perim=18.46u w=4.615u l=4.615u
XR2 iovss sub / ptap1 r=208.667m A=4.43n Perim=266.24u w=66.56u l=66.56u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Corner
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Corner iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XR1 vss sub / ptap1 r=35.383 A=13.177p Perim=14.52u w=3.63u l=3.63u
XR0 iovss sub / ptap1 r=93.041m A=10.13n Perim=402.6u w=100.65u l=100.65u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Filler400
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Filler400 iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XR1 vss sub / ptap1 r=246.192 A=680.625f Perim=3.3u w=825n l=825n
XR0 iovss sub / ptap1 r=6.246 A=114.169p Perim=42.74u w=10.685u l=10.685u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Filler200
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Filler200 iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XR1 vss sub / ptap1 r=246.192 A=680.625f Perim=3.3u w=825n l=825n
XR0 iovss sub / ptap1 r=14.724 A=40.96p Perim=25.6u w=6.4u l=6.4u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Filler1000
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Filler1000 iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XR1 vss sub / ptap1 r=162.013 A=1.369p Perim=4.68u w=1.17u l=1.17u
XR0 iovss sub / ptap1 r=2.443 A=328.697p Perim=72.52u w=18.13u l=18.13u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Filler2000
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Filler2000 iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XR1 vss sub / ptap1 r=101.912 A=2.856p Perim=6.76u w=1.69u l=1.69u
XR0 iovss sub / ptap1 r=1.224 A=695.113p Perim=105.46u w=26.365u l=26.365u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Filler10000
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Filler10000 iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XR1 vss sub / ptap1 r=32.364 A=14.861p Perim=15.42u w=3.855u l=3.855u
XR0 iovss sub / ptap1 r=253.731m A=3.622n Perim=240.72u w=60.18u l=60.18u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_P20N0D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_P20N0D iovdd iovss pad sub
*.PININFO iovdd:B iovss:B pad:B
MP0 pad net2 iovdd iovdd sg13_hv_pmos m=1 w=266.4u l=600.0n ng=40
*RR0 net2 iovdd 6.768K $SUB=iovdd $[res_rppd] m=1 l=12.9u w=500n ps=180n 
+ trise=0.0 b=0
RR0 iovdd net2 rppd m=1 l=12.9u w=500n
+ trise=0.0 b=0
XR1 iovss sub / ptap1 r=9.826 A=66.994p Perim=32.74u w=8.185u l=8.185u
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_Clamp_N20N0D
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_Clamp_N20N0D iovss pad sub
*.PININFO iovss:B pad:B
MN0 pad net2 iovss sub sg13_hv_nmos m=1 w=88.000u l=600.0n ng=20
XR0 iovss sub / ptap1 r=11.438 A=55.801p Perim=29.88u w=7.47u l=7.47u
*RR1 iovss net2 1.959K $SUB=sub $[res_rppd] m=1 l=3.54u w=500n ps=180n 
+ trise=0.0 b=0
RR1 iovss net2 rppd m=1 l=3.54u w=500n
+ trise=0.0 b=0
.ENDS

************************************************************************
* Library Name: sg13g2_io
* Cell Name:    sg13g2_IOPadAnalog
* View Name:    schematic
************************************************************************

.SUBCKT sg13g2_IOPadAnalog iovdd iovss pad padres vdd vss sub
*.PININFO iovdd:B iovss:B pad:B padres:B vdd:B vss:B
XI9 iovdd iovss pad sub / sg13g2_Clamp_P20N0D
XI3 iovss pad iovdd sub / sg13g2_DCNDiode
XI2 pad iovdd iovss sub / sg13g2_DCPDiode
*** WHYYYYYY. Lets put it like that for now. My god this is annoying
*XI6 padres iovss pad iovdda sub / sg13g2_SecondaryProtection
XI6 padres iovss pad iovdd sub / sg13g2_SecondaryProtection
XI8 iovss pad sub / sg13g2_Clamp_N20N0D
XR1 vss sub / ptap1 r=22.579 A=23.863p Perim=19.54u w=4.885u l=4.885u
XR2 iovss sub / ptap1 r=214.8m A=4.3n Perim=262.3u w=65.575u l=65.575u
.ENDS
.SUBCKT sg13g2_bpd60
.ENDS

.SUBCKT sg13g2_bpd70
.ENDS

.SUBCKT sg13g2_bpd80
.ENDS
*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

.SUBCKT sg13g2_Clamp_N20N0DExt iovss pad sub
*.PININFO iovss:B pad:B
MN0 pad net2 iovss sub sg13_hv_nmos m=1 w=88.000u l=600.0n ng=20
XR0 iovss sub / ptap1 r=11.438 A=55.801p Perim=29.88u w=7.47u l=7.47u
*RR1 iovss net2 1.959K $SUB=sub $[res_rppd] m=1 l=3.54u w=500n ps=180n 
+ trise=0.0 b=0
*RR0 net2 iovdd 6.768K $SUB=iovdd $[res_rppd] m=1 l=12.9u w=500n ps=180n 
+ trise=0.0 b=0
RR0 iovdd net2 rppd m=1 l=12.9u w=500n
+ trise=0.0 b=0
.ENDS

.SUBCKT sg13g2_SecondaryProtectionExt core minus pad plus sub
*.PININFO core:B minus:B pad:B plus:B
*RR0 pad core 586.899 $SUB=sub $[res_rppd] m=1 l=2u w=1u ps=180n trise=0.0 b=0
RR0 pad core rppd m=1 l=2u w=1u
DD0 sub core dantenna m=1 w=640n l=3.1u a=1.984p p=7.48u
XR1 minus sub / ptap1 r=46.556 A=9.03p Perim=12.02u w=3.005u l=3.005u
DD1 core plus dpantenna m=1 w=640n l=4.98u a=3.187p p=11.24u
.ENDS

.SUBCKT sg13g2_Clamp_P20N0DExt iovdd iovss pad sub
*.PININFO iovdd:B iovss:B pad:B
MP0 pad net2 iovdd iovdd sg13_hv_pmos m=1 w=266.4u l=600.0n ng=40
RR0 net2 iovdd 6.768K $SUB=iovdd $[res_rppd] m=1 l=12.9u w=500n ps=180n 
+ trise=0.0 b=0
XR1 iovss sub / ptap1 r=9.826 A=66.994p Perim=32.74u w=8.185u l=8.185u
.ENDS

.SUBCKT sg13g2_RCClampInverterExt in iovss out supply sub
*.PININFO in:B iovss:B out:B supply:B
MN1 iovss in iovss sub sg13_hv_nmos m=1 w=126.000u l=9.5u ng=14
MN0 out in iovss sub sg13_hv_nmos m=1 w=108.000u l=500.0n ng=12
XR0 iovss sub / ptap1 r=9.59 A=68.973p Perim=33.22u w=8.305u l=8.305u
MP0 out in supply supply sg13_hv_pmos m=1 w=350.000u l=500.0n ng=50
.ENDS

.SUBCKT sg13g2_RCClampResistorExt pin1 pin2 sub
*.PININFO pin1:B pin2:B
R$274 pin2 pin1 rppd w=1u l=520u ps=0 b=0 m=1
.ENDS

.SUBCKT sg13g2_RCClampResistorExt_Orig pin1 pin2 sub
*.PININFO pin1:B pin2:B
RR29 net15 net16 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR28 net20 net21 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR27 net23 net24 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR24 net17 net18 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR23 net16 net17 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR21 net25 pin2 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR20 net22 net23 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR19 net19 net20 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR17 net24 net25 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR16 net21 net22 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR15 net18 net19 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR14 net5 net6 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR13 net8 net9 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR12 net11 net12 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR11 net14 net15 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR10 net2 net3 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR9 net1 net2 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR8 net13 net14 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR7 net10 net11 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR6 net7 net8 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR5 net4 net5 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR4 net12 net13 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR3 net9 net10 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 
+ b=0
RR2 net6 net7 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR1 net3 net4 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
RR0 pin1 net1 5.239K $SUB=sub $[res_rppd] m=1 l=20u w=1u ps=180n trise=0.0 b=0
.ENDS

.SUBCKT sg13g2_Clamp_N43N43D4RExt gate pad tie sub
*.PININFO gate:I pad:B tie:B
MN0<1> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<2> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<3> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<4> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<5> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<6> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<7> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<8> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<9> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<10> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<11> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<12> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<13> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<14> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<15> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<16> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<17> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<18> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<19> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<20> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<21> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<22> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<23> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<24> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<25> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<26> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<27> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<28> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<29> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<30> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<31> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<32> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<33> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<34> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<35> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<36> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<37> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<38> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<39> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<40> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<41> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<42> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<43> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<44> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<45> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<46> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<47> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<48> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<49> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<50> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<51> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<52> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<53> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<54> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<55> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<56> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<57> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<58> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<59> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<60> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<61> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<62> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<63> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<64> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<65> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<66> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<67> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<68> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<69> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<70> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<71> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<72> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<73> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<74> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<75> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<76> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<77> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<78> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<79> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<80> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<81> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<82> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<83> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<84> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<85> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<86> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<87> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<88> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<89> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<90> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<91> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<92> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<93> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<94> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<95> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<96> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<97> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<98> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<99> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<100> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<101> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<102> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<103> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<104> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<105> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<106> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<107> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<108> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<109> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<110> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<111> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<112> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<113> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<114> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<115> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<116> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<117> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<118> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<119> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<120> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<121> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<122> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<123> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<124> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<125> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<126> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<127> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<128> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<129> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<130> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<131> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<132> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<133> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<134> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<135> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<136> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<137> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<138> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<139> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<140> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<141> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<142> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<143> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<144> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<145> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<146> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<147> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<148> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<149> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<150> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<151> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<152> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<153> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<154> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<155> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<156> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<157> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<158> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<159> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<160> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<161> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<162> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<163> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<164> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<165> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<166> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<167> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<168> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<169> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<170> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<171> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
MN0<172> pad gate tie sub sg13_hv_nmos m=1 w=4.4u l=600.0n ng=1
XR0 tie sub / ptap1 r=9.999 A=65.61p Perim=32.4u w=8.1u l=8.1u
DD0 sub gate dantenna m=1 w=480n l=480n a=230.4f p=1.92u
.ENDS

.SUBCKT sg13g2_DCNDiodeExt anode cathode guard sub
*.PININFO anode:B cathode:B guard:B
DD1 sub cathode dantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
DD0 sub cathode dantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
XR0 anode sub / ptap1 r=5.191 A=141.253p Perim=47.54u w=11.885u l=11.885u
.ENDS

.SUBCKT sg13g2_DCPDiodeExt anode cathode guard sub
*.PININFO anode:B cathode:B guard:B
DD1 anode cathode dpantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
DD0 anode cathode dpantenna m=1 w=1.26u l=27.78u a=35.003p p=58.08u
XR0 guard sub / ptap1 r=17.289 A=33.524p Perim=23.16u w=5.79u l=5.79u
.ENDS

.SUBCKT sg13g2_IOPadVssExt iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
XI1 iovss vss iovss sub / sg13g2_DCNDiodeExt
XI2 vss iovdd iovss sub / sg13g2_DCPDiodeExt
XR1 iovss sub / ptap1 r=174.346m A=5.329n Perim=292u w=73u l=73u
XR0 vss sub / ptap1 r=22.832 A=23.523p Perim=19.4u w=4.85u l=4.85u
.ENDS

.SUBCKT sg13g2_IOPadVddExt iovdd iovss vdd vss sub
*.PININFO iovdd:B iovss:B vdd:B vss:B
* OHH MY GOD
*XI0 net2 vdd iovssa sub / sg13g2_Clamp_N43N43D4RExt
XI0 net2 vdd iovss sub / sg13g2_Clamp_N43N43D4RExt
XI2 vdd net1 sub / sg13g2_RCClampResistorExt
XR1 iovss sub / ptap1 r=456.33m A=1.97n Perim=177.54u w=44.385u l=44.385u
XR0 vss sub / ptap1 r=22.472 A=24.01p Perim=19.6u w=4.9u l=4.9u
XI1 net1 iovss net2 vdd sub  / sg13g2_RCClampInverterExt
.ENDS

.SUBCKT sg13g2_IOPadAVDD iovdd iovss pad padres vdd vss sub
*.PININFO iovdd:B iovss:B pad:B padres:B vdd:B vss:B
XI9 iovdd iovss pad sub / sg13g2_Clamp_P20N0DExt
XI3 iovss pad iovdd sub / sg13g2_DCNDiodeExt
XI2 pad iovdd iovss sub / sg13g2_DCPDiodeExt
XI6 padres iovss pad iovdd sub / sg13g2_SecondaryProtectionExt
XI8 iovss pad sub / sg13g2_Clamp_N20N0DExt
XR1 vss sub / ptap1 r=22.579 A=23.863p Perim=19.54u w=4.885u l=4.885u
XR2 iovss sub / ptap1 r=214.8m A=4.3n Perim=262.3u w=65.575u l=65.575u
.ENDS
.SUBCKT sealring
.ENDS
** Created by: circuit_gen.AN2D0
** Cell name: AN2D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_AN2D0 a1 a2 vdd vss z
*.PININFO a1:B a2:B vdd:B vss:B z:B 
M_u2_M_u3 net6 a1 x_u2_net6 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u3_M_u2 z net6 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u2_M_u4 x_u2_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u3_M_u3 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u2_M_u2 net6 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u2_M_u1 net6 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.AN2D1
** Cell name: AN2D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_AN2D1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
M_u2_M_u3 net6 a1 x_u2_net6 vss sg13_lv_nmos l=1.300e-07 w=6.550e-07
M_u3_M_u2 z net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_M_u4 x_u2_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.550e-07
M_u3_M_u3 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_M_u2 net6 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_M_u1 net6 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.AN2D2
** Cell name: AN2D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_AN2D2 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
M_u2_M_u3 net10 a1 x_u2_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_M_u2_0 z net10 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_M_u2_1 z net10 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_M_u4 x_u2_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_M_u3_0 z net10 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_M_u3_1 z net10 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_M_u2 net10 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_M_u1 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.AN2D4
** Cell name: AN2D4
** Lib name: sg13g2f
.SUBCKT sg13g2f_AN2D4 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
M_u2_0_M_u3 p0 a1 x_u2_0_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_0_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_1_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_2_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_3_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_0_M_u4 x_u2_0_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_1_M_u4 x_u2_1_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_1_M_u3 p0 a1 x_u2_1_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_0_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_1_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_2_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_3_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_0_M_u2 p0 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_0_M_u1 p0 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_1_M_u2 p0 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_1_M_u1 p0 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.AO21D0
** Cell name: AO21D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_AO21D0 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI7 net32 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7 net59 a1 net32 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI6 net59 b vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI8_M_u2 z net59 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u3 net22 a1 net59 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI8_M_u3 z net59 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u4 net22 a2 net59 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u2 net22 b vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.AO21D1
** Cell name: AO21D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_AO21D1 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI7 net32 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u7 net59 a1 net32 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI6 net59 b vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI8_M_u2 z net59 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3 net22 a1 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI8_M_u3 z net59 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u4 net22 a2 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2 net22 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.AO21D2
** Cell name: AO21D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_AO21D2 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI7 net32 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u7 net59 a1 net32 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI6 net59 b vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI8_0_M_u2 z net59 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI8_1_M_u2 z net59 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3 net22 a1 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI8_0_M_u3 z net59 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI8_1_M_u3 z net59 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u4 net22 a2 net59 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2 net22 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.AOI21D0
** Cell name: AOI21D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_AOI21D0 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
MI2 zn a1 net27 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI7 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI6 zn b vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI5 zn a2 net13 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u2 net13 b vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI4 zn a1 net13 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.AOI21D1
** Cell name: AOI21D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_AOI21D1 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
MI2 zn a1 net27 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI3 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u7 zn b vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u4 net13 a2 zn vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2 net13 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3 net13 a1 zn vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.ANTENNA
** Cell name: ANTENNA
** Lib name: sg13g2f
.SUBCKT sg13g2f_ANTENNA i vdd vss
*.PININFO i:I vdd:B vss:B
Ddn_1 vss i dantenna m=1 w=1.485u l=970n a=1440.45f
DD0 i vdd dpantenna m=1 w=1.485u l=970n a=1440.45f
.ENDS

** Created by: circuit_gen.BUFFD0
** Cell name: BUFFD0
** Lib name: sg13g2f
.SUBCKT sg13g2f_BUFFD0 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u3_M_u2 z net6 vss vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
M_u2_M_u2 net6 i vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07
M_u3_M_u3 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=5.850e-07
M_u2_M_u3 net6 i vdd vdd sg13_lv_pmos l=1.300e-07 w=3.600e-07
.ENDS

** Created by: circuit_gen.BUFFD1
** Cell name: BUFFD1
** Lib name: sg13g2f
.SUBCKT sg13g2f_BUFFD1 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u3_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_M_u2 net8 i vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u3_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_M_u3 net8 i vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.BUFFD2
** Cell name: BUFFD2
** Lib name: sg13g2f
.SUBCKT sg13g2f_BUFFD2 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u2_M_u2 net8 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_0_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_1_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_M_u3 net8 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_0_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_1_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.BUFFD4
** Cell name: BUFFD4
** Lib name: sg13g2f
.SUBCKT sg13g2f_BUFFD4 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u3_0_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_1_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_2_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_3_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_0_M_u2 p0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2_1_M_u2 p0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3_0_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_1_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_2_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u3_3_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_0_M_u3 p0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2_1_M_u3 p0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.BUFFD6
** Cell name: BUFFD6
** Lib name: sg13g2f
.SUBCKT sg13g2f_BUFFD6 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u2_M_u2_0 net8 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=1
M_u2_M_u2_1 net8 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=0
M_u3_0_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=1
M_u3_1_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=0
M_u3_2_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=1
M_u3_3_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=0
M_u3_4_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=1
M_u3_5_M_u2 z net8 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=0
M_u2_M_u3_0 net8 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=1
M_u2_M_u3_1 net8 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=0
M_u3_0_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=1
M_u3_1_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=0
M_u3_2_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=1
M_u3_3_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=0
M_u3_4_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=1
M_u3_5_M_u3 z net8 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=0
.ENDS

** Created by: circuit_gen.BUFFD8
** Cell name: BUFFD8
** Lib name: sg13g2f
.SUBCKT sg13g2f_BUFFD8 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
MI1_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=0
MI2_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=4.850e-07 $pos=1 $flip=1
M_u2_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=0
M_u7_0_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=1
M_u7_1_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=0
M_u7_2_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=1
M_u7_3_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=0
M_u7_4_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=1
M_u7_5_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=8 $flip=0
M_u7_6_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=9 $flip=1
M_u7_7_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=10 $flip=0
MI1_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=0
MI2_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=8.050e-07 $pos=1 $flip=1
M_u2_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
M_u7_0_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=1
M_u7_1_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=0
M_u7_2_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
M_u7_3_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
M_u7_4_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=1
M_u7_5_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=8 $flip=0
M_u7_6_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=1
M_u7_7_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=0
.ENDS

** Created by: circuit_gen.BUFFD12
** Cell name: BUFFD12
** Lib name: sg13g2f
.SUBCKT sg13g2f_BUFFD12 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
M_u2_0_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=4.300e-07 $pos=0 $flip=0
M_u2_1_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=4.300e-07 $pos=1 $flip=1
M_u2_2_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=4.300e-07 $pos=2 $flip=0
M_u2_3_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=4.300e-07 $pos=3 $flip=1
M_u2_4_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=4.300e-07 $pos=4 $flip=0
MU8_0_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=1
MU8_1_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=0
MU8_2_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=1
MU8_3_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=8 $flip=0
MU8_4_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=9 $flip=1
MU8_5_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=10 $flip=0
MU8_6_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=11 $flip=1
MU8_7_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=12 $flip=0
MU8_8_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=13 $flip=1
MU8_9_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=14 $flip=0
MU8_10_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=15 $flip=1
MU8_11_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=16 $flip=0
M_u2_0_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=0
M_u2_1_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=1
M_u2_2_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=0
M_u2_3_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=1
M_u2_4_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=0
MU8_0_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
MU8_1_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
MU8_2_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=1
MU8_3_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=8 $flip=0
MU8_4_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=1
MU8_5_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=0
MU8_6_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=11 $flip=1
MU8_7_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=12 $flip=0
MU8_8_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=13 $flip=1
MU8_9_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=14 $flip=0
MU8_10_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=15 $flip=1
MU8_11_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=16 $flip=0
.ENDS

** Created by: circuit_gen.BUFFD16
** Cell name: BUFFD16
** Lib name: sg13g2f
.SUBCKT sg13g2f_BUFFD16 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
MI6_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=2.500e-07 $pos=0 $flip=1
M_u2_0_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=0
M_u2_1_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=1
M_u2_2_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=0
M_u2_3_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=1
M_u2_4_M_u2 n0 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=0
MU8_0_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=1
MU8_1_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=0
MU8_2_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=8 $flip=1
MU8_3_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=9 $flip=0
MU8_4_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=10 $flip=1
MU8_5_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=11 $flip=0
MU8_6_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=12 $flip=1
MU8_7_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=13 $flip=0
MU8_8_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=14 $flip=1
MU8_9_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=15 $flip=0
MU8_10_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=16 $flip=1
MU8_11_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=17 $flip=0
MU8_12_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=18 $flip=1
MU8_13_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=19 $flip=0
MU8_14_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=20 $flip=1
MU8_15_M_u2 z n0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=21 $flip=0
MI6_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=3.950e-07 $pos=0 $flip=1
M_u2_0_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=0
M_u2_1_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=1
M_u2_2_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=0
M_u2_3_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=1
M_u2_4_M_u3 n0 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=0
MU8_0_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=1
MU8_1_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=0
MU8_2_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=8 $flip=1
MU8_3_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=0
MU8_4_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=1
MU8_5_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=11 $flip=0
MU8_6_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=12 $flip=1
MU8_7_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=13 $flip=0
MU8_8_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=14 $flip=1
MU8_9_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=15 $flip=0
MU8_10_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=16 $flip=1
MU8_11_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=17 $flip=0
MU8_12_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=18 $flip=1
MU8_13_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=19 $flip=0
MU8_14_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=20 $flip=1
MU8_15_M_u3 z n0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=21 $flip=0
.ENDS

** Created by: circuit_gen.DEL0
** Cell name: DEL0
** Lib name: sg13g2f
.SUBCKT sg13g2f_DEL0 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
MI2_M_u2 z net3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU7_M_u2 net3 net5 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU5_M_u2 net5 net9 vss vss sg13_lv_nmos l=1.300e-07 w=4.800e-07
MI1_M_u2 net9 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI2_M_u3 z net3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU7_M_u3 net3 net5 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.040e-06
MU5_M_u3 net5 net9 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u3 net9 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.DEL2
** Cell name: DEL2
** Lib name: sg13g2f
.SUBCKT sg13g2f_DEL2 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
MI2_M_u2 z net3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU7_M_u2 net3 net5 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU5_M_u2 net5 net9 vss vss sg13_lv_nmos l=1.300e-07 w=4.800e-07
MI1_M_u2 net9 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI2_M_u3 z net3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU7_M_u3 net3 net5 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.000e-07
MU5_M_u3 net5 net9 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u3 net9 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.DEL02
** Cell name: DEL02
** Lib name: sg13g2f
.SUBCKT sg13g2f_DEL02 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
MI17 net3 net21 net27 vss sg13_lv_nmos l=1.300e-07 w=3.350e-07
MI18 net27 net21 vss vss sg13_lv_nmos l=1.300e-07 w=3.350e-07
MI5 net21 net9 net24 vss sg13_lv_nmos l=1.300e-07 w=3.350e-07
MI16 net24 net9 vss vss sg13_lv_nmos l=1.300e-07 w=3.350e-07
MI2_M_u2 z net3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u2 net9 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI15 net27 net21 net3 vdd sg13_lv_pmos l=1.300e-07 w=5.650e-07
MI13 net24 net9 net21 vdd sg13_lv_pmos l=1.300e-07 w=5.650e-07
MI3 vdd net9 net24 vdd sg13_lv_pmos l=1.300e-07 w=5.650e-07
MI14 vdd net21 net27 vdd sg13_lv_pmos l=1.300e-07 w=5.650e-07
MI2_M_u3 z net3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u3 net9 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.DEL4
** Cell name: DEL4
** Lib name: sg13g2f
.SUBCKT sg13g2f_DEL4 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
MI2_M_u2 z net13 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU7_M_u2 net13 net11 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU5_M_u2 net11 net9 vss vss sg13_lv_nmos l=1.300e-07 w=4.800e-07
MI1_M_u2 net9 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI2_M_u3 z net13 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU7_M_u3 net13 net11 vdd vdd sg13_lv_pmos l=1.300e-07 w=8.500e-07
MU5_M_u3 net11 net9 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u3 net9 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.DEL005
** Cell name: DEL005
** Lib name: sg13g2f
.SUBCKT sg13g2f_DEL005 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
MI12 net3 i net22 vss sg13_lv_nmos l=1.300e-07 w=4.250e-07
MI13 net22 i vss vss sg13_lv_nmos l=1.300e-07 w=4.250e-07
MI2_M_u2 z net3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI10 net3 i net21 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI3 net21 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI2_M_u3 z net3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.DEL015
** Cell name: DEL015
** Lib name: sg13g2f
.SUBCKT sg13g2f_DEL015 i vdd vss z
*.PININFO i:I z:O vdd:B vss:B 
MI11 net27 net21 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI10 net3 net21 net27 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI5 net21 net9 net24 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI111 net24 net9 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI2_M_u2 z net3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u2 net9 i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI8 net27 net21 net3 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI9 vdd net21 net27 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI4 net24 net9 net21 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI3 vdd net9 net24 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI2_M_u3 z net3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u3 net9 i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.DFCNQD1
** Cell name: DFCNQD1
** Lib name: sg13g2
.SUBCKT sg13g2f_DFCNQD1 cdn cp d q vdd vss
*.PININFO cdn:I cp:I d:I q:O vdd:B vss:B 
Mcpbn incpb cp vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07 $pos=0 $flip=0
Mcpbp incpb cp vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07 $pos=0 $flip=0
Mcpn incp incpb vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07 $pos=1 $flip=1
Mcpp incp incpb vdd vdd sg13_lv_pmos l=1.300e-07 w=5.500e-07 $pos=1 $flip=1
MI4 net52 incpb vss vss sg13_lv_nmos l=1.300e-07 w=3.500e-07 $pos=3 $flip=1
MI7 net85 incp vdd vdd sg13_lv_pmos l=1.300e-07 w=8.100e-07 $pos=3 $flip=1
Mdd0n d0 d net52 vss sg13_lv_nmos l=1.300e-07 w=3.500e-07 $pos=4 $flip=1
Mdd0p d0 d net85 vdd sg13_lv_pmos l=1.300e-07 w=8.100e-07 $pos=4 $flip=1
MI47 d0 incp net59 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=5 $flip=0
MI45 d0 incpb net98 vdd sg13_lv_pmos l=1.300e-07 w=3.300e-07 $pos=5 $flip=0
MI48 net59 d1 net62 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=6 $flip=0
MI43 net98 d1 vdd vdd sg13_lv_pmos l=1.300e-07 w=3.050e-07 $pos=6 $flip=0
Mcdn0n net62 cdn vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=7 $flip=0
Md0d1n d1 d0 vss vss sg13_lv_nmos l=1.300e-07 w=4.300e-07 $pos=8 $flip=1
Mcdn0p net98 cdn vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07 $pos=8 $flip=0
Mswd1d2n d1 incp d2 vss sg13_lv_nmos l=1.300e-07 w=4.900e-07 $pos=9 $flip=0
Mdod1p d1 d0 vdd vdd sg13_lv_pmos l=1.300e-07 w=7.150e-07 $pos=9 $flip=1
MI23 d2 incpb net57 vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=10 $flip=0
Mswd1d2p d1 incpb d2 vdd sg13_lv_pmos l=1.300e-07 w=1.030e-06 $pos=10 $flip=0
MI26 d2 incp net88 vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07 $pos=11 $flip=0
MI24 net57 d3 vss vss sg13_lv_nmos l=1.300e-07 w=2.450e-07 $pos=12 $flip=0
MI28 net88 d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=2.750e-07 $pos=12 $flip=0
Mcdn1n net37 cdn vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07 $pos=13 $flip=1
Mcdn1p d3 cdn vdd vdd sg13_lv_pmos l=1.300e-07 w=9.900e-07 $pos=13 $flip=1
Md2d3n d3 d2 net37 vss sg13_lv_nmos l=1.300e-07 w=7.000e-07 $pos=14 $flip=1
Md2d3p d3 d2 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.900e-07 $pos=14 $flip=0
Mobp q d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.100e-06 $pos=15 $flip=1
Mobn q d3 vss vss sg13_lv_nmos l=1.300e-07 w=7.000e-07 $pos=16 $flip=1
.ENDS

** Created by: circuit_gen.DFQD1
** Cell name: DFQD1
** Lib name: sg13g2f
.SUBCKT sg13g2f_DFQD1 cp d q vdd vss
*.PININFO cp:I d:I q:O vdd:B vss:B 
MI4 net43 incpb vss vss sg13_lv_nmos l=1.300e-07 w=4.200e-07
MI23 d2 incpb net42 vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI5 d0 d net43 vss sg13_lv_nmos l=1.300e-07 w=4.200e-07
MI47 d0 incp net50 vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI48 net50 d1 vss vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI24 net42 d3 vss vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI50 d1 incp d2 vss sg13_lv_nmos l=1.300e-07 w=3.850e-07
MI32_M_u2 incp incpb vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI31_M_u2 incpb cp vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI27_M_u2 q d3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI53_M_u2 d3 d2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI13_M_u2 d1 d0 vss vss sg13_lv_nmos l=1.300e-07 w=4.700e-07
MI6 d0 d net66 vdd sg13_lv_pmos l=1.300e-07 w=7.500e-07
MI32_M_u3 incp incpb vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI31_M_u3 incpb cp vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI27_M_u3 q d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI53_M_u3 d3 d2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI13_M_u3 d1 d0 vdd vdd sg13_lv_pmos l=1.300e-07 w=7.500e-07
MI7 net66 incp vdd vdd sg13_lv_pmos l=1.300e-07 w=8.850e-07
MI52 d1 incpb d2 vdd sg13_lv_pmos l=1.300e-07 w=1.065e-06
MI28 net74 d3 vdd vdd sg13_lv_pmos l=1.300e-07 w=3.000e-07
MI26 d2 incp net74 vdd sg13_lv_pmos l=1.300e-07 w=3.000e-07
MI45 d0 incpb net84 vdd sg13_lv_pmos l=1.300e-07 w=3.000e-07
MI43 net84 d1 vdd vdd sg13_lv_pmos l=1.300e-07 w=3.000e-07
.ENDS

** Created by: circuit_gen.FILL1
** Cell name: FILL1
** Lib name: sg13g2f
.SUBCKT sg13g2f_FILL1 vdd vss
*.PININFO vdd:B vss:B 
.ENDS

** Created by: circuit_gen.FILL2
** Cell name: FILL2
** Lib name: sg13g2f
.SUBCKT sg13g2f_FILL2 vdd vss
*.PININFO vdd:B vss:B 
.ENDS

** Created by: circuit_gen.FILL4
** Cell name: FILL4
** Lib name: sg13g2f
.SUBCKT sg13g2f_FILL4 vdd vss
*.PININFO vdd:B vss:B 
.ENDS

** Created by: circuit_gen.FILL8
** Cell name: FILL8
** Lib name: sg13g2f
.SUBCKT sg13g2f_FILL8 vdd vss
*.PININFO vdd:B vss:B 
.ENDS

** Created by: circuit_gen.INVD0
** Cell name: INVD0
** Lib name: sg13g2f
.SUBCKT sg13g2f_INVD0 i vdd vss zn
*.PININFO i:I zn:O vdd:B vss:B 
MU1_M_u2 zn i vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU1_M_u3 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.INVD1
** Cell name: INVD1
** Lib name: sg13g2f
.SUBCKT sg13g2f_INVD1 i z vss vdd
*.PININFO i:I z:O vss:B vdd:B
M0 z i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M1 z i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.INVD2
** Cell name: INVD2
** Lib name: sg13g2f
.SUBCKT sg13g2f_INVD2 i vdd vss zn
*.PININFO i:I zn:O vdd:B vss:B 
MU1_M_u2_0 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_M_u2_1 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_M_u3_0 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_M_u3_1 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.INVD4
** Cell name: INVD4
** Lib name: sg13g2f
.SUBCKT sg13g2f_INVD4 i vdd vss zn
*.PININFO i:I zn:O vdd:B vss:B 
MU1_M_u2_0 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_M_u2_1 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_M_u2_2 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_M_u2_3 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_M_u3_0 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_M_u3_1 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_M_u3_2 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_M_u3_3 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.INVD6
** Cell name: INVD6
** Lib name: sg13g2f
.SUBCKT sg13g2f_INVD6 i vdd vss zn
*.PININFO i:I zn:O vdd:B vss:B 
MU1_M_u2_0 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=0
MU1_M_u2_1 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=1
MU1_M_u2_2 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=0
MU1_M_u2_3 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=1
MU1_M_u2_4 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=0
MU1_M_u2_5 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=1
MU1_M_u3_0 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=0
MU1_M_u3_1 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MU1_M_u3_2 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
MU1_M_u3_3 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=1
MU1_M_u3_4 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=0
MU1_M_u3_5 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
.ENDS

** Created by: circuit_gen.INVD8
** Cell name: INVD8
** Lib name: sg13g2f
.SUBCKT sg13g2f_INVD8 i vdd vss zn
*.PININFO i:I zn:O vdd:B vss:B 
MU1_M_u2_0 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=0
MU1_M_u2_1 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=1
MU1_M_u2_2 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=0
MU1_M_u2_3 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=1
MU1_M_u2_4 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=0
MU1_M_u2_5 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=1
MU1_M_u2_6 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=0
MU1_M_u2_7 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=1
MU1_M_u3_0 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=0
MU1_M_u3_1 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MU1_M_u3_2 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
MU1_M_u3_3 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=1
MU1_M_u3_4 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=0
MU1_M_u3_5 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
MU1_M_u3_6 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
MU1_M_u3_7 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=1
.ENDS

** Created by: circuit_gen.INVD12
** Cell name: INVD12
** Lib name: sg13g2f
.SUBCKT sg13g2f_INVD12 i vdd vss zn
*.PININFO i:I zn:O vdd:B vss:B 
MU1_M_u2_0 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=0
MU1_M_u2_1 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=1
MU1_M_u2_2 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=0
MU1_M_u2_3 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=1
MU1_M_u2_4 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=0
MU1_M_u2_5 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=1
MU1_M_u2_6 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=0
MU1_M_u2_7 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=1
MU1_M_u2_8 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=8 $flip=0
MU1_M_u2_9 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=9 $flip=1
MU1_M_u2_10 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=10 $flip=0
MU1_M_u2_11 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=11 $flip=1
MU1_M_u3_0 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=0
MU1_M_u3_1 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MU1_M_u3_2 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
MU1_M_u3_3 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=1
MU1_M_u3_4 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=0
MU1_M_u3_5 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
MU1_M_u3_6 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
MU1_M_u3_7 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=1
MU1_M_u3_8 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=8 $flip=0
MU1_M_u3_9 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=1
MU1_M_u3_10 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=0
MU1_M_u3_11 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=11 $flip=1
.ENDS

** Created by: circuit_gen.INVD16
** Cell name: INVD16
** Lib name: sg13g2f
.SUBCKT sg13g2f_INVD16 i vdd vss zn
*.PININFO i:I zn:O vdd:B vss:B 
MU1_M_u2_0 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=0
MU1_M_u2_1 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=1
MU1_M_u2_2 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=0
MU1_M_u2_3 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=1
MU1_M_u2_4 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=0
MU1_M_u2_5 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=1
MU1_M_u2_6 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=0
MU1_M_u2_7 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=1
MU1_M_u2_8 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=8 $flip=0
MU1_M_u2_9 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=9 $flip=1
MU1_M_u2_10 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=10 $flip=0
MU1_M_u2_11 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=11 $flip=1
MU1_M_u2_12 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=12 $flip=0
MU1_M_u2_13 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=13 $flip=1
MU1_M_u2_14 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=14 $flip=0
MU1_M_u2_15 zn i vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=15 $flip=1
MU1_M_u3_0 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=0
MU1_M_u3_1 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MU1_M_u3_2 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
MU1_M_u3_3 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=1
MU1_M_u3_4 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=0
MU1_M_u3_5 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
MU1_M_u3_6 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
MU1_M_u3_7 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=1
MU1_M_u3_8 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=8 $flip=0
MU1_M_u3_9 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=1
MU1_M_u3_10 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=0
MU1_M_u3_11 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=11 $flip=1
MU1_M_u3_12 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=12 $flip=0
MU1_M_u3_13 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=13 $flip=1
MU1_M_u3_14 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=14 $flip=0
MU1_M_u3_15 zn i vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=15 $flip=1
.ENDS

** Created by: circuit_gen.MUX2D0
** Cell name: MUX2D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_MUX2D0 i0 i1 s vdd vss z
*.PININFO i0:I i1:I s:I z:O vdd:B vss:B 
MI15_M_u3 net46 s net28 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU7_M_u3 net48 net42 net28 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI16_M_u2 net48 i0 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI17_M_u2 net46 i1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI18_M_u2 net42 s vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU29_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI15_M_u2 net46 net42 net28 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MU7_M_u2 net48 s net28 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI16_M_u3 net48 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI17_M_u3 net46 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI18_M_u3 net42 s vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MU29_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.MUX2D1
** Cell name: MUX2D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_MUX2D1 i0 i1 s vdd vss z
*.PININFO i0:I i1:I s:I z:O vdd:B vss:B 
MI15_M_u3 net46 s net28 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU7_M_u3 net48 net42 net28 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI20_M_u2 net46 i1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI19_M_u2 net48 i0 vss vss sg13_lv_nmos l=1.300e-07 w=5.200e-07
MI18_M_u2 net42 s vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU29_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI15_M_u2 net46 net42 net28 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MU7_M_u2 net48 s net28 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI20_M_u3 net46 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI19_M_u3 net48 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.900e-07
MI18_M_u3 net42 s vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MU29_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=8.400e-07
.ENDS

** Created by: circuit_gen.MUX2D2
** Cell name: MUX2D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_MUX2D2 i0 i1 s vdd vss z
*.PININFO i0:I i1:I s:I z:O vdd:B vss:B 
MI15_M_u3 net46 s net28 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU7_M_u3 net48 net42 net28 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI20_M_u2 net46 i1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI19_M_u2 net48 i0 vss vss sg13_lv_nmos l=1.300e-07 w=5.200e-07
MI18_M_u2 net42 s vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU29_0_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU29_1_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI15_M_u2 net46 net42 net28 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MU7_M_u2 net48 s net28 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI20_M_u3 net46 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI19_M_u3 net48 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.900e-07
MI18_M_u3 net42 s vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MU29_0_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU29_1_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.MUX2D4
** Cell name: MUX2D4
** Lib name: sg13g2f
.SUBCKT sg13g2f_MUX2D4 i0 i1 s vdd vss z
*.PININFO i0:I i1:I s:I z:O vdd:B vss:B 
MI21_M_u3 net24 s net28 vss sg13_lv_nmos l=1.300e-07 w=6.200e-07
MU7_M_u3 net16 net42 net28 vss sg13_lv_nmos l=1.300e-07 w=5.350e-07
MI20_0_M_u2 net24 i1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI20_1_M_u2 net24 i1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI19_0_M_u2 net16 i0 vss vss sg13_lv_nmos l=1.300e-07 w=5.200e-07
MI19_1_M_u2 net16 i0 vss vss sg13_lv_nmos l=1.300e-07 w=5.200e-07
MI18_M_u2 net42 s vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU29_0_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU29_1_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU29_2_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU29_3_M_u2 z net28 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI21_M_u2 net24 net42 net28 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU7_M_u2 net16 s net28 vdd sg13_lv_pmos l=1.300e-07 w=1.095e-06
MI20_0_M_u3 net24 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI20_1_M_u3 net24 i1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI19_0_M_u3 net16 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.750e-07
MI19_1_M_u3 net16 i0 vdd vdd sg13_lv_pmos l=1.300e-07 w=9.750e-07
MI18_M_u3 net42 s vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MU29_0_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU29_1_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU29_2_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU29_3_M_u3 z net28 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.ND2D0
** Cell name: ND2D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_ND2D0 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI0_M_u3 zn a1 xi0_net6 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI0_M_u4 xi0_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI0_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI0_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.ND2D1
** Cell name: ND2D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_ND2D1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u3 zn a1 xi1_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u4 xi1_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.ND2D2
** Cell name: ND2D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_ND2D2 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MU3_0_M_u3 zn a1 xu3_0_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU3_0_M_u4 xu3_0_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU3_1_M_u4 xu3_1_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU3_1_M_u3 zn a1 xu3_1_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU3_0_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU3_0_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU3_1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU3_1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.ND2D4
** Cell name: ND2D4
** Lib name: sg13g2f
.SUBCKT sg13g2f_ND2D4 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_0_M_u3 zn a1 xi1_0_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_0_M_u4 xi1_0_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_1_M_u4 xi1_1_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_1_M_u3 zn a1 xi1_1_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_2_M_u4 xi1_2_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_2_M_u3 zn a1 xi1_2_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_3_M_u4 xi1_3_net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_3_M_u3 zn a1 xi1_3_net6 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_0_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_0_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_2_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_2_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_3_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_3_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.ND3D0
** Cell name: ND3D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_ND3D0 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
MI2_M_u4 zn a1 xi2_net10 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI2_M_u5 xi2_net10 a2 xi2_net13 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI2_M_u6 xi2_net13 a3 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI2_M_u3 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI2_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI2_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.ND3D1
** Cell name: ND3D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_ND3D1 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 xi1_net10 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u5 xi1_net10 a2 xi1_net13 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u6 xi1_net13 a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u3 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.ND3D2
** Cell name: ND3D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_ND3D2 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
MI0_0_M_u4 zn a1 xi0_0_net10 vss sg13_lv_nmos l=1.300e-07 w=6.700e-07
MI0_0_M_u5 xi0_0_net10 a2 xi0_0_net13 vss sg13_lv_nmos l=1.300e-07 w=6.700e-07
MI0_0_M_u6 xi0_0_net13 a3 vss vss sg13_lv_nmos l=1.300e-07 w=6.700e-07
MI0_1_M_u4 zn a1 xi0_1_net10 vss sg13_lv_nmos l=1.300e-07 w=6.700e-07
MI0_1_M_u5 xi0_1_net10 a2 xi0_1_net13 vss sg13_lv_nmos l=1.300e-07 w=6.700e-07
MI0_1_M_u6 xi0_1_net13 a3 vss vss sg13_lv_nmos l=1.300e-07 w=6.700e-07
MI0_0_M_u3 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI0_0_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI0_0_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI0_1_M_u3 zn a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI0_1_M_u1 zn a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI0_1_M_u2 zn a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.NR2D0
** Cell name: NR2D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_NR2D0 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI1_M_u3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI1_M_u2 zn a1 xi1_net8 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI1_M_u1 xi1_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.NR2D1
** Cell name: NR2D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_NR2D1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_M_u4 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1_M_u2 zn a1 xi1_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1_M_u1 xi1_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.NR2D2
** Cell name: NR2D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_NR2D2 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI1_0_M_u3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=1
MI1_0_M_u4 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=0
MI1_1_M_u4 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=1
MI1_1_M_u3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=0
MI1_0_M_u1 xi1_0_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=1
MI1_0_M_u2 zn a1 xi1_0_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MI1_1_M_u2 zn a1 xi1_1_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
MI1_1_M_u1 xi1_1_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=0
.ENDS

** Created by: circuit_gen.NR2D4
** Cell name: NR2D4
** Lib name: sg13g2f
.SUBCKT sg13g2f_NR2D4 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI6_0 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=1
MI15_0 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=0
MI15_1 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=1
MI6_2 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=0
MI6_3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=1
MI15_2 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=0
MI15_3 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=1
MI6_1 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=0
MI27_0 net26_0_ a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=1
MI28_0 zn a1 net26_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MI28_1 zn a1 net26_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
MI27_1 net26_1_ a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=0
MI27_2 net26_2_ a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=1
MI28_2 zn a1 net26_2_ vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
MI28_3 zn a1 net26_3_ vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
MI27_3 net26_3_ a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=0
.ENDS

** Created by: circuit_gen.NR3D0
** Cell name: NR3D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_NR3D0 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
M_u4 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI2 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI3 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI0 net28 a2 net25 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u1 net25 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI1 zn a1 net28 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.NR3D1
** Cell name: NR3D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_NR3D1 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
M_u4 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=1
MI2 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=0
MI3 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=1
M_u1_0 net34_0_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=1
MI4_0 net37_0_ a2 net34_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MI5_0 zn a1 net37_0_ vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=1
MI5_1 zn a1 net37_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=0
MI4_1 net37_1_ a2 net34_1_ vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=0
M_u1_1 net34_1_ a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=0
.ENDS

** Created by: circuit_gen.NR3D2
** Cell name: NR3D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_NR3D2 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
M_u4_0 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=1
M_u4_1 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=0
MI6_0 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=1
MI6_1 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=0
MI7_0 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=9 $flip=1
MI7_1 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=10 $flip=0
M_u1_0 net34 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=0
M_u1_1 net34 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
M_u1_2 net34 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
M_u1_3 net34 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=1
MI22_0 net31 a2 net34 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=1
MI22_1 net31 a2 net34 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=0
MI22_2 net31 a2 net34 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=1
MI22_3 net31 a2 net34 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=0
MI23_0 zn a1 net31 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=1
MI23_1 zn a1 net31 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=0
MI23_2 zn a1 net31 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=11 $flip=1
MI23_3 zn a1 net31 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=12 $flip=0
.ENDS

** Created by: circuit_gen.NR3D4
** Cell name: NR3D4
** Lib name: sg13g2f
.SUBCKT sg13g2f_NR3D4 a1 a2 a3 vdd vss zn
*.PININFO a1:I a2:I a3:I zn:O vdd:B vss:B 
MI0_M_u4_0 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=1
MI0_M_u4_1 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=0
MI0_M_u4_2 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=1
MI0_M_u4_3 zn a3 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=0
MI0_M_u5_0 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=12 $flip=1
MI0_M_u5_1 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=13 $flip=0
MI0_M_u5_2 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=14 $flip=1
MI0_M_u5_3 zn a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=15 $flip=0
MI0_M_u6_0 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=17 $flip=1
MI0_M_u6_1 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=18 $flip=0
MI0_M_u6_2 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=19 $flip=1
MI0_M_u6_3 zn a1 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=20 $flip=0
MI0_M_u1_0 xi0_net9 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=0
MI0_M_u1_1 xi0_net9 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MI0_M_u1_2 xi0_net9 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
MI0_M_u1_3 xi0_net9 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=1
MI0_M_u1_4 xi0_net9 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=0
MI0_M_u1_5 xi0_net9 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
MI0_M_u1_6 xi0_net9 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
MI0_M_u1_7 xi0_net9 a3 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=1
MI0_M_u2_0 xi0_net12 a2 xi0_net9 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=8 $flip=1
MI0_M_u2_1 xi0_net12 a2 xi0_net9 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=0
MI0_M_u2_2 xi0_net12 a2 xi0_net9 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=1
MI0_M_u2_3 xi0_net12 a2 xi0_net9 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=11 $flip=0
MI0_M_u2_4 xi0_net12 a2 xi0_net9 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=12 $flip=1
MI0_M_u2_5 xi0_net12 a2 xi0_net9 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=13 $flip=0
MI0_M_u2_6 xi0_net12 a2 xi0_net9 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=14 $flip=1
MI0_M_u2_7 xi0_net12 a2 xi0_net9 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=15 $flip=0
MI0_M_u3_0 zn a1 xi0_net12 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=17 $flip=1
MI0_M_u3_1 zn a1 xi0_net12 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=18 $flip=0
MI0_M_u3_2 zn a1 xi0_net12 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=19 $flip=1
MI0_M_u3_3 zn a1 xi0_net12 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=20 $flip=0
MI0_M_u3_4 zn a1 xi0_net12 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=21 $flip=1
MI0_M_u3_5 zn a1 xi0_net12 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=22 $flip=0
MI0_M_u3_6 zn a1 xi0_net12 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=23 $flip=1
MI0_M_u3_7 zn a1 xi0_net12 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=24 $flip=0
.ENDS

** Created by: circuit_gen.OA21D1
** Cell name: OA21D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_OA21D1 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI12 net14 a2 net20 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI11 net14 a1 net20 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI6 net20 b vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI8_M_u2 z net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI9 net14 a1 net24 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI8_M_u3 z net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2 net14 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI7 net24 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.OA21D2
** Cell name: OA21D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_OA21D2 a1 a2 b vdd vss z
*.PININFO a1:I a2:I b:I z:O vdd:B vss:B 
MI12 net14 a2 net20 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI11 net14 a1 net20 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI6 net20 b vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI8_0_M_u2 z net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI8_1_M_u2 z net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI9 net14 a1 net24 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI8_0_M_u3 z net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI8_1_M_u3 z net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u2 net14 b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI7 net24 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.OAI21D0
** Cell name: OAI21D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_OAI21D0 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
M_u2 zn a1 net15 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u3 zn a2 net15 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u4 net15 b vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI16_MI12 zn a1 xi16_net11 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u9 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI16_MI13 xi16_net11 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.OAI21D1
** Cell name: OAI21D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_OAI21D1 a1 a2 b vdd vss zn
*.PININFO a1:I a2:I b:I zn:O vdd:B vss:B 
M_u2 zn a1 net15 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3 zn a2 net15 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u4 net15 b vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI16_MI12 zn a1 xi16_net11 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u9 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI16_MI13 xi16_net11 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.OAI211D0
** Cell name: OAI211D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_OAI211D0 a1 a2 b c vdd vss zn
*.PININFO a1:I a2:I b:I c:I zn:O vdd:B vss:B 
MI8 net36 b net24 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI9 net24 c vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u2 zn a1 net36 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI7 zn a2 net36 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI6 zn a2 net35 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI5 net35 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI4 zn c vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u12 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.OAI211D1
** Cell name: OAI211D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_OAI211D1 a1 a2 b c vdd vss zn
*.PININFO a1:I a2:I b:I c:I zn:O vdd:B vss:B 
MI2 net36 b net24 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI3 net24 c vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u2 zn a1 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u3 zn a2 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI1 zn a2 net35 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI0 net35 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u11 zn c vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u12 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.OAI211D4
** Cell name: OAI211D4
** Lib name: sg13g2f
.SUBCKT sg13g2f_OAI211D4 a1 a2 b c vdd vss zn
*.PININFO a1:I a2:I b:I c:I zn:O vdd:B vss:B 
MI13_0 zn a2 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=0
MI13_1 zn a2 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=1
MI13_2 zn a2 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=0
MI13_3 zn a2 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=1
MI14_0 zn a1 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=0
MI14_1 zn a1 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=1
MI14_2 zn a1 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=0
MI14_3 zn a1 net36 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=1
MI2_0 net36 b net24 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=9 $flip=1
MI2_1 net36 b net24 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=10 $flip=0
MI2_2 net36 b net24 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=11 $flip=1
MI2_3 net36 b net24 vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=12 $flip=0
MI12_0 net24 c vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=13 $flip=0
MI12_1 net24 c vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=14 $flip=1
MI12_2 net24 c vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=15 $flip=0
MI12_3 net24 c vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=16 $flip=1
MI11_0 zn a2 net35 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=1
MI11_1 zn a2 net35 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=0
MI11_2 zn a2 net35 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=1
MI11_3 zn a2 net35 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=0
MI9_0 net35 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
MI9_1 net35 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
MI9_2 net35 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=1
MI9_3 net35 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=8 $flip=0
M_u12_0 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=1
M_u12_1 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=0
M_u12_2 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=11 $flip=1
M_u12_3 zn b vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=12 $flip=0
MI8_0 zn c vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=13 $flip=1
MI8_1 zn c vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=14 $flip=0
MI8_2 zn c vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=15 $flip=1
MI8_3 zn c vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=16 $flip=0
.ENDS

** Created by: circuit_gen.OR2D0
** Cell name: OR2D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_OR2D0 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MU1_M_u2 z net7 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_M_u4 net7 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_M_u3 net7 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_M_u2 net7 a1 x_u7_net8 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MU1_M_u3 z net7 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u7_M_u1 x_u7_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.OR2D1
** Cell name: OR2D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_OR2D1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MU1_M_u2 z net7 vss vss sg13_lv_nmos l=1.300e-07 w=6.550e-07
M_u7_M_u4 net7 a1 vss vss sg13_lv_nmos l=1.300e-07 w=6.550e-07
M_u7_M_u3 net7 a2 vss vss sg13_lv_nmos l=1.300e-07 w=6.550e-07
M_u7_M_u2 net7 a1 x_u7_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_M_u3 z net7 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u7_M_u1 x_u7_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.OR2D2
** Cell name: OR2D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_OR2D2 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MU1_0_M_u2 z net9 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_1_M_u2 z net9 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u7_M_u4 net9 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_M_u3 net9 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_M_u2 net9 a1 x_u7_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_0_M_u3 z net9 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_1_M_u3 z net9 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u7_M_u1 x_u7_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.OR2D4
** Cell name: OR2D4
** Lib name: sg13g2f
.SUBCKT sg13g2f_OR2D4 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MU1_0_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_1_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_2_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MU1_3_M_u2 z p0 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u7_0_M_u4 p0 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_0_M_u3 p0 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_1_M_u4 p0 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_1_M_u3 p0 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_0_M_u2 p0 a1 x_u7_0_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_0_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_1_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_2_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MU1_3_M_u3 z p0 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u7_0_M_u1 x_u7_0_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u7_1_M_u1 x_u7_1_net8 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u7_1_M_u2 p0 a1 x_u7_1_net8 vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.TAPCELL
** Cell name: TAPCELL
** Lib name: sg13g2f
.SUBCKT sg13g2f_TAPCELL vdd vss
*.PININFO vdd:B vss:B 
.ENDS

** Created by: circuit_gen.TIEH
** Cell name: TIEH
** Lib name: sg13g2f
.SUBCKT sg13g2f_TIEH vdd vss z
*.PININFO z:O vdd:B vss:B 
M_u2 net6 net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u1 z net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.TIEL
** Cell name: TIEL
** Lib name: sg13g2f
.SUBCKT sg13g2f_TIEL vdd vss zn
*.PININFO zn:O vdd:B vss:B 
M_u2 zn net6 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u1 net6 net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
.ENDS

** Created by: circuit_gen.XNR2D0
** Cell name: XNR2D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_XNR2D0 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
MI2_M_u3 net28 net10 net14 vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI0_M_u3 net6 a1 net14 vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI1_M_u2 net28 net6 vss vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
M_u2_M_u2 net6 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u4_M_u2 zn net14 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u8_M_u2 net10 a1 vss vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI2_M_u2 net28 a1 net14 vdd sg13_lv_pmos l=1.300e-07 w=4.050e-07
MI0_M_u2 net6 net10 net14 vdd sg13_lv_pmos l=1.300e-07 w=4.050e-07
MI1_M_u3 net28 net6 vdd vdd sg13_lv_pmos l=1.300e-07 w=4.050e-07
M_u2_M_u3 net6 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u4_M_u3 zn net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u8_M_u3 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=4.050e-07
.ENDS

** Created by: circuit_gen.XNR2D1
** Cell name: XNR2D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_XNR2D1 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
M_u2_M_u2 net4 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u5_M_u2 net6 net4 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u4_M_u2 zn net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u8_M_u2 net10 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u6_M_u3 net4 a1 net14 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_M_u3 net6 net10 net14 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u6_M_u2 net4 net10 net14 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u2_M_u3 net4 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u5_M_u3 net6 net4 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u4_M_u3 zn net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u8_M_u3 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u7_M_u2 net6 a1 net14 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.XNR2D2
** Cell name: XNR2D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_XNR2D2 a1 a2 vdd vss zn
*.PININFO a1:I a2:I zn:O vdd:B vss:B 
M_u6_M_u3 net4 a1 net14 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u7_M_u3 net6 net10 net14 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u2_M_u2 net4 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u5_M_u2 net6 net4 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u4_0_M_u2 zn net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u4_1_M_u2 zn net14 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
M_u8_M_u2 net10 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u6_M_u2 net4 net10 net14 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u7_M_u2 net6 a1 net14 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u2_M_u3 net4 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u5_M_u3 net6 net4 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u4_0_M_u3 zn net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u4_1_M_u3 zn net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
M_u8_M_u3 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.XOR2D0
** Cell name: XOR2D0
** Lib name: sg13g2f
.SUBCKT sg13g2f_XOR2D0 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MI5_M_u3 net25 a1 net14 vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
M_u6_M_u3 net4 net10 net14 vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI6_M_u2 net25 net4 vss vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI1_M_u2 net4 a2 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
M_u4_M_u2 z net14 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI2_M_u2 net10 a1 vss vss sg13_lv_nmos l=1.300e-07 w=2.500e-07
MI5_M_u2 net25 net10 net14 vdd sg13_lv_pmos l=1.300e-07 w=4.050e-07
M_u6_M_u2 net4 a1 net14 vdd sg13_lv_pmos l=1.300e-07 w=4.050e-07
MI6_M_u3 net25 net4 vdd vdd sg13_lv_pmos l=1.300e-07 w=4.050e-07
MI1_M_u3 net4 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
M_u4_M_u3 z net14 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI2_M_u3 net10 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=4.050e-07
.ENDS

** Created by: circuit_gen.XOR2D1
** Cell name: XOR2D1
** Lib name: sg13g2f
.SUBCKT sg13g2f_XOR2D1 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MI6_M_u3 net41 a1 net21 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI2_M_u3 net27 net23 net21 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI7_M_u2 net41 net27 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI3_M_u2 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI4_M_u2 z net21 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI5_M_u2 net23 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI6_M_u2 net41 net23 net21 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI2_M_u2 net27 a1 net21 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI7_M_u3 net41 net27 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI3_M_u3 net27 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI4_M_u3 z net21 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI5_M_u3 net23 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS

** Created by: circuit_gen.XOR2D2
** Cell name: XOR2D2
** Lib name: sg13g2f
.SUBCKT sg13g2f_XOR2D2 a1 a2 vdd vss z
*.PININFO a1:I a2:I z:O vdd:B vss:B 
MI6_M_u3 net41 a1 net21 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI2_M_u3 net27 net23 net21 vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI7_M_u2 net41 net27 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI3_M_u2 net27 a2 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI4_0_M_u2 z net21 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI4_1_M_u2 z net21 vss vss sg13_lv_nmos l=1.300e-07 w=7.200e-07
MI5_M_u2 net23 a1 vss vss sg13_lv_nmos l=1.300e-07 w=3.600e-07
MI6_M_u2 net41 net23 net21 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI2_M_u2 net27 a1 net21 vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI7_M_u3 net41 net27 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
MI3_M_u3 net27 a2 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI4_0_M_u3 z net21 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI4_1_M_u3 z net21 vdd vdd sg13_lv_pmos l=1.300e-07 w=1.200e-06
MI5_M_u3 net23 a1 vdd vdd sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS
** Cell name: SARADC_CELL_INVX0_ASSW
** Lib name: sg13g2f
.SUBCKT SARADC_CELL_INVX0_ASSW i vdd vss zn vnw vpw
*.PININFO i:B zn:B vdd:B vss:B 
MU1_M_u2 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=3.600e-07
MU1_M_u3 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=6.000e-07
.ENDS
** Cell name: SARADC_CELL_INVX16_ASCAP
** Lib name: sg13g2f
.SUBCKT SARADC_CELL_INVX16_ASCAP i vdd vss zn vnw vpw
*.PININFO i:I zn:O vdd:B vss:B 
MU1_M_u2_0 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=0 $flip=0
MU1_M_u2_1 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=1 $flip=1
MU1_M_u2_2 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=2 $flip=0
MU1_M_u2_3 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=3 $flip=1
MU1_M_u2_4 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=4 $flip=0
MU1_M_u2_5 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=5 $flip=1
MU1_M_u2_6 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=6 $flip=0
MU1_M_u2_7 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=7 $flip=1
MU1_M_u2_8 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=8 $flip=0
MU1_M_u2_9 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=9 $flip=1
MU1_M_u2_10 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=10 $flip=0
MU1_M_u2_11 zn i vss vpw sg13_lv_nmos l=1.300e-07 w=7.200e-07 $pos=11 $flip=1
MU1_M_u3_0 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=0 $flip=0
MU1_M_u3_1 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=1 $flip=1
MU1_M_u3_2 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=2 $flip=0
MU1_M_u3_3 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=3 $flip=1
MU1_M_u3_4 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=4 $flip=0
MU1_M_u3_5 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=5 $flip=1
MU1_M_u3_6 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=6 $flip=0
MU1_M_u3_7 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=7 $flip=1
MU1_M_u3_8 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=8 $flip=0
MU1_M_u3_9 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=9 $flip=1
MU1_M_u3_10 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=10 $flip=0
MU1_M_u3_11 zn i vdd vnw sg13_lv_pmos l=1.300e-07 w=1.200e-06 $pos=11 $flip=1
.ENDS
** Cell name: SARADC_FILLTIE2
** Lib name: sg13g2f
.SUBCKT SARADC_FILLTIE2 vdd vss
*.PININFO vdd:B vss:B 
.ENDS
** Cell name: SARADC_FILL1
.SUBCKT SARADC_FILL1 vdd vss
*.PININFO vdd:B vss:B 
.ENDS
** Cell name: SARADC_FILL1_NOPOWER
.SUBCKT SARADC_FILL1_NOPOWER
.ENDS
* CDL Netlist generated by OpenROAD

*.BUSDELIMITER [

.SUBCKT SARADC AVDD CLK GO RESULT[0] RESULT[1] RESULT[2] RESULT[3]
+ RESULT[4] RST SAMPLE VALID VDD VIN VIP VREFH VREFL VSS
Xanalog/buflogic.conv.cmpbegin.ccmpbuf1.impl analog/buflogic.conv.cmpbegin.CCMPNR
+ AVDD VSS analog/buflogic.conv.cmpbegin.CCMPNR1 sg13g2f_BUFFD8
Xanalog/buflogic.conv.cmpbegin.ccmpbuf2.impl analog/buflogic.conv.cmpbegin.CCMPNR1
+ AVDD VSS analog/buflogic.CMP sg13g2f_BUFFD16
Xanalog/buflogic.conv.cmpbegin.ccmpnor.impl SAMPLE CLKBUF
+ VALID AVDD VSS analog/buflogic.conv.cmpbegin.CCMPNR sg13g2f_NR3D4
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.ibuf16.impl RESULTN\[1\]
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZL sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.ln1.impl analog/buflogic.conv.re2cr\[1\].ren2crh.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZNL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.ln2.impl analog/buflogic.conv.re2cr\[1\].ren2crh.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zbuf.impl analog/buflogic.conv.re2cr\[1\].ren2crh.ZLD3
+ AVDD VSS analog/CRH\[0\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zdel_1.impl1 analog/buflogic.conv.re2cr\[1\].ren2crh.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.zdel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zdel_1.impl2 analog/buflogic.conv.re2cr\[1\].ren2crh.zdel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zdel_2.impl1 analog/buflogic.conv.re2cr\[1\].ren2crh.ZLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.zdel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zdel_2.impl2 analog/buflogic.conv.re2cr\[1\].ren2crh.zdel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zdel_3.impl1 analog/buflogic.conv.re2cr\[1\].ren2crh.ZLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.zdel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zdel_3.impl2 analog/buflogic.conv.re2cr\[1\].ren2crh.zdel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.znbuf.impl analog/buflogic.conv.re2cr\[1\].ren2crh.ZNLD3
+ AVDD VSS analog/CRHB\[0\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zndel_1.impl1 analog/buflogic.conv.re2cr\[1\].ren2crh.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.zndel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zndel_1.impl2 analog/buflogic.conv.re2cr\[1\].ren2crh.zndel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZNLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zndel_2.impl1 analog/buflogic.conv.re2cr\[1\].ren2crh.ZNLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.zndel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zndel_2.impl2 analog/buflogic.conv.re2cr\[1\].ren2crh.zndel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZNLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zndel_3.impl1 analog/buflogic.conv.re2cr\[1\].ren2crh.ZNLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.zndel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].ren2crh.zndel_3.impl2 analog/buflogic.conv.re2cr\[1\].ren2crh.zndel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].ren2crh.ZNLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.ibuf16.impl RESULT[1]
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZL sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.ln1.impl analog/buflogic.conv.re2cr\[1\].rep2crl.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZNL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.ln2.impl analog/buflogic.conv.re2cr\[1\].rep2crl.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zbuf.impl analog/buflogic.conv.re2cr\[1\].rep2crl.ZLD3
+ AVDD VSS analog/CRL\[0\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zdel_1.impl1 analog/buflogic.conv.re2cr\[1\].rep2crl.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.zdel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zdel_1.impl2 analog/buflogic.conv.re2cr\[1\].rep2crl.zdel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zdel_2.impl1 analog/buflogic.conv.re2cr\[1\].rep2crl.ZLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.zdel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zdel_2.impl2 analog/buflogic.conv.re2cr\[1\].rep2crl.zdel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zdel_3.impl1 analog/buflogic.conv.re2cr\[1\].rep2crl.ZLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.zdel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zdel_3.impl2 analog/buflogic.conv.re2cr\[1\].rep2crl.zdel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.znbuf.impl analog/buflogic.conv.re2cr\[1\].rep2crl.ZNLD3
+ AVDD VSS analog/CRLB\[0\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zndel_1.impl1 analog/buflogic.conv.re2cr\[1\].rep2crl.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.zndel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zndel_1.impl2 analog/buflogic.conv.re2cr\[1\].rep2crl.zndel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZNLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zndel_2.impl1 analog/buflogic.conv.re2cr\[1\].rep2crl.ZNLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.zndel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zndel_2.impl2 analog/buflogic.conv.re2cr\[1\].rep2crl.zndel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZNLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zndel_3.impl1 analog/buflogic.conv.re2cr\[1\].rep2crl.ZNLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.zndel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[1\].rep2crl.zndel_3.impl2 analog/buflogic.conv.re2cr\[1\].rep2crl.zndel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[1\].rep2crl.ZNLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.ibuf16.impl RESULTN\[2\]
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZL sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.ln1.impl analog/buflogic.conv.re2cr\[2\].ren2crh.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZNL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.ln2.impl analog/buflogic.conv.re2cr\[2\].ren2crh.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zbuf.impl analog/buflogic.conv.re2cr\[2\].ren2crh.ZLD3
+ AVDD VSS analog/CRH\[1\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zdel_1.impl1 analog/buflogic.conv.re2cr\[2\].ren2crh.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.zdel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zdel_1.impl2 analog/buflogic.conv.re2cr\[2\].ren2crh.zdel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zdel_2.impl1 analog/buflogic.conv.re2cr\[2\].ren2crh.ZLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.zdel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zdel_2.impl2 analog/buflogic.conv.re2cr\[2\].ren2crh.zdel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zdel_3.impl1 analog/buflogic.conv.re2cr\[2\].ren2crh.ZLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.zdel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zdel_3.impl2 analog/buflogic.conv.re2cr\[2\].ren2crh.zdel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.znbuf.impl analog/buflogic.conv.re2cr\[2\].ren2crh.ZNLD3
+ AVDD VSS analog/CRHB\[1\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zndel_1.impl1 analog/buflogic.conv.re2cr\[2\].ren2crh.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.zndel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zndel_1.impl2 analog/buflogic.conv.re2cr\[2\].ren2crh.zndel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZNLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zndel_2.impl1 analog/buflogic.conv.re2cr\[2\].ren2crh.ZNLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.zndel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zndel_2.impl2 analog/buflogic.conv.re2cr\[2\].ren2crh.zndel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZNLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zndel_3.impl1 analog/buflogic.conv.re2cr\[2\].ren2crh.ZNLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.zndel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].ren2crh.zndel_3.impl2 analog/buflogic.conv.re2cr\[2\].ren2crh.zndel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].ren2crh.ZNLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.ibuf16.impl RESULT[2]
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZL sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.ln1.impl analog/buflogic.conv.re2cr\[2\].rep2crl.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZNL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.ln2.impl analog/buflogic.conv.re2cr\[2\].rep2crl.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zbuf.impl analog/buflogic.conv.re2cr\[2\].rep2crl.ZLD3
+ AVDD VSS analog/CRL\[1\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zdel_1.impl1 analog/buflogic.conv.re2cr\[2\].rep2crl.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.zdel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zdel_1.impl2 analog/buflogic.conv.re2cr\[2\].rep2crl.zdel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zdel_2.impl1 analog/buflogic.conv.re2cr\[2\].rep2crl.ZLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.zdel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zdel_2.impl2 analog/buflogic.conv.re2cr\[2\].rep2crl.zdel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zdel_3.impl1 analog/buflogic.conv.re2cr\[2\].rep2crl.ZLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.zdel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zdel_3.impl2 analog/buflogic.conv.re2cr\[2\].rep2crl.zdel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.znbuf.impl analog/buflogic.conv.re2cr\[2\].rep2crl.ZNLD3
+ AVDD VSS analog/CRLB\[1\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zndel_1.impl1 analog/buflogic.conv.re2cr\[2\].rep2crl.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.zndel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zndel_1.impl2 analog/buflogic.conv.re2cr\[2\].rep2crl.zndel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZNLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zndel_2.impl1 analog/buflogic.conv.re2cr\[2\].rep2crl.ZNLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.zndel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zndel_2.impl2 analog/buflogic.conv.re2cr\[2\].rep2crl.zndel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZNLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zndel_3.impl1 analog/buflogic.conv.re2cr\[2\].rep2crl.ZNLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.zndel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[2\].rep2crl.zndel_3.impl2 analog/buflogic.conv.re2cr\[2\].rep2crl.zndel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[2\].rep2crl.ZNLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.ibuf16.impl RESULTN\[3\]
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZL sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.ln1.impl analog/buflogic.conv.re2cr\[3\].ren2crh.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZNL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.ln2.impl analog/buflogic.conv.re2cr\[3\].ren2crh.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zbuf.impl analog/buflogic.conv.re2cr\[3\].ren2crh.ZLD3
+ AVDD VSS analog/CRH\[2\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zdel_1.impl1 analog/buflogic.conv.re2cr\[3\].ren2crh.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.zdel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zdel_1.impl2 analog/buflogic.conv.re2cr\[3\].ren2crh.zdel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zdel_2.impl1 analog/buflogic.conv.re2cr\[3\].ren2crh.ZLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.zdel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zdel_2.impl2 analog/buflogic.conv.re2cr\[3\].ren2crh.zdel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zdel_3.impl1 analog/buflogic.conv.re2cr\[3\].ren2crh.ZLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.zdel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zdel_3.impl2 analog/buflogic.conv.re2cr\[3\].ren2crh.zdel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.znbuf.impl analog/buflogic.conv.re2cr\[3\].ren2crh.ZNLD3
+ AVDD VSS analog/CRHB\[2\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zndel_1.impl1 analog/buflogic.conv.re2cr\[3\].ren2crh.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.zndel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zndel_1.impl2 analog/buflogic.conv.re2cr\[3\].ren2crh.zndel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZNLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zndel_2.impl1 analog/buflogic.conv.re2cr\[3\].ren2crh.ZNLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.zndel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zndel_2.impl2 analog/buflogic.conv.re2cr\[3\].ren2crh.zndel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZNLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zndel_3.impl1 analog/buflogic.conv.re2cr\[3\].ren2crh.ZNLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.zndel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].ren2crh.zndel_3.impl2 analog/buflogic.conv.re2cr\[3\].ren2crh.zndel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].ren2crh.ZNLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.ibuf16.impl RESULT[3]
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZL sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.ln1.impl analog/buflogic.conv.re2cr\[3\].rep2crl.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZNL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.ln2.impl analog/buflogic.conv.re2cr\[3\].rep2crl.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zbuf.impl analog/buflogic.conv.re2cr\[3\].rep2crl.ZLD3
+ AVDD VSS analog/CRL\[2\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zdel_1.impl1 analog/buflogic.conv.re2cr\[3\].rep2crl.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.zdel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zdel_1.impl2 analog/buflogic.conv.re2cr\[3\].rep2crl.zdel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zdel_2.impl1 analog/buflogic.conv.re2cr\[3\].rep2crl.ZLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.zdel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zdel_2.impl2 analog/buflogic.conv.re2cr\[3\].rep2crl.zdel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zdel_3.impl1 analog/buflogic.conv.re2cr\[3\].rep2crl.ZLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.zdel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zdel_3.impl2 analog/buflogic.conv.re2cr\[3\].rep2crl.zdel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.znbuf.impl analog/buflogic.conv.re2cr\[3\].rep2crl.ZNLD3
+ AVDD VSS analog/CRLB\[2\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zndel_1.impl1 analog/buflogic.conv.re2cr\[3\].rep2crl.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.zndel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zndel_1.impl2 analog/buflogic.conv.re2cr\[3\].rep2crl.zndel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZNLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zndel_2.impl1 analog/buflogic.conv.re2cr\[3\].rep2crl.ZNLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.zndel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zndel_2.impl2 analog/buflogic.conv.re2cr\[3\].rep2crl.zndel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZNLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zndel_3.impl1 analog/buflogic.conv.re2cr\[3\].rep2crl.ZNLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.zndel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[3\].rep2crl.zndel_3.impl2 analog/buflogic.conv.re2cr\[3\].rep2crl.zndel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[3\].rep2crl.ZNLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.ibuf16.impl RESULTN\[4\]
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZL sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.ln1.impl analog/buflogic.conv.re2cr\[4\].ren2crh.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZNL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.ln2.impl analog/buflogic.conv.re2cr\[4\].ren2crh.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zbuf.impl analog/buflogic.conv.re2cr\[4\].ren2crh.ZLD3
+ AVDD VSS analog/CRH\[3\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zdel_1.impl1 analog/buflogic.conv.re2cr\[4\].ren2crh.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.zdel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zdel_1.impl2 analog/buflogic.conv.re2cr\[4\].ren2crh.zdel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zdel_2.impl1 analog/buflogic.conv.re2cr\[4\].ren2crh.ZLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.zdel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zdel_2.impl2 analog/buflogic.conv.re2cr\[4\].ren2crh.zdel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zdel_3.impl1 analog/buflogic.conv.re2cr\[4\].ren2crh.ZLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.zdel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zdel_3.impl2 analog/buflogic.conv.re2cr\[4\].ren2crh.zdel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.znbuf.impl analog/buflogic.conv.re2cr\[4\].ren2crh.ZNLD3
+ AVDD VSS analog/CRHB\[3\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zndel_1.impl1 analog/buflogic.conv.re2cr\[4\].ren2crh.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.zndel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zndel_1.impl2 analog/buflogic.conv.re2cr\[4\].ren2crh.zndel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZNLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zndel_2.impl1 analog/buflogic.conv.re2cr\[4\].ren2crh.ZNLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.zndel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zndel_2.impl2 analog/buflogic.conv.re2cr\[4\].ren2crh.zndel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZNLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zndel_3.impl1 analog/buflogic.conv.re2cr\[4\].ren2crh.ZNLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.zndel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].ren2crh.zndel_3.impl2 analog/buflogic.conv.re2cr\[4\].ren2crh.zndel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].ren2crh.ZNLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.ibuf16.impl RESULT[4]
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZL sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.ln1.impl analog/buflogic.conv.re2cr\[4\].rep2crl.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZNL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.ln2.impl analog/buflogic.conv.re2cr\[4\].rep2crl.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZL sg13g2f_INVD8
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zbuf.impl analog/buflogic.conv.re2cr\[4\].rep2crl.ZLD3
+ AVDD VSS analog/CRL\[3\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zdel_1.impl1 analog/buflogic.conv.re2cr\[4\].rep2crl.ZL
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.zdel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zdel_1.impl2 analog/buflogic.conv.re2cr\[4\].rep2crl.zdel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zdel_2.impl1 analog/buflogic.conv.re2cr\[4\].rep2crl.ZLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.zdel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zdel_2.impl2 analog/buflogic.conv.re2cr\[4\].rep2crl.zdel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zdel_3.impl1 analog/buflogic.conv.re2cr\[4\].rep2crl.ZLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.zdel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zdel_3.impl2 analog/buflogic.conv.re2cr\[4\].rep2crl.zdel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.znbuf.impl analog/buflogic.conv.re2cr\[4\].rep2crl.ZNLD3
+ AVDD VSS analog/CRLB\[3\] sg13g2f_BUFFD16
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zndel_1.impl1 analog/buflogic.conv.re2cr\[4\].rep2crl.ZNL
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.zndel_1.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zndel_1.impl2 analog/buflogic.conv.re2cr\[4\].rep2crl.zndel_1.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZNLD1 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zndel_2.impl1 analog/buflogic.conv.re2cr\[4\].rep2crl.ZNLD1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.zndel_2.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zndel_2.impl2 analog/buflogic.conv.re2cr\[4\].rep2crl.zndel_2.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZNLD2 sg13g2f_BUFFD2
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zndel_3.impl1 analog/buflogic.conv.re2cr\[4\].rep2crl.ZNLD2
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.zndel_3.Z1
+ sg13g2f_DEL4
Xanalog/buflogic.conv.re2cr\[4\].rep2crl.zndel_3.impl2 analog/buflogic.conv.re2cr\[4\].rep2crl.zndel_3.Z1
+ AVDD VSS analog/buflogic.conv.re2cr\[4\].rep2crl.ZNLD3 sg13g2f_BUFFD2
Xanalog/buflogic.conv.smpcs.choldb.impl analog/buflogic.HOLD
+ AVDD VSS analog/buflogic.conv.smpcs.CHOLDB sg13g2f_INVD8
Xanalog/buflogic.conv.smpcs.choldb1.impl analog/buflogic.conv.smpcs.CHOLDB
+ AVDD VSS analog/buflogic.conv.smpcs.CHOLDB1 sg13g2f_BUFFD8
Xanalog/buflogic.conv.smpcs.clkbuf.impl clknet_1_0__leaf_CLK_regs
+ AVDD VSS CLKBUF sg13g2f_BUFFD16
Xanalog/buflogic.conv.smpcs.clkbufd1.impl1 CLKBUF AVDD VSS
+ analog/buflogic.conv.smpcs.clkbufd1.Z1 sg13g2f_DEL4
Xanalog/buflogic.conv.smpcs.clkbufd1.impl2 analog/buflogic.conv.smpcs.clkbufd1.Z1
+ AVDD VSS analog/buflogic.conv.smpcs.CLKBUFD1 sg13g2f_BUFFD4
Xanalog/buflogic.conv.smpcs.clkbufd2.impl1 analog/buflogic.conv.smpcs.CLKBUFD1
+ AVDD VSS analog/buflogic.conv.smpcs.clkbufd2.Z1 sg13g2f_DEL4
Xanalog/buflogic.conv.smpcs.clkbufd2.impl2 analog/buflogic.conv.smpcs.clkbufd2.Z1
+ AVDD VSS analog/buflogic.conv.smpcs.CLKBUFD2 sg13g2f_BUFFD4
Xanalog/buflogic.conv.smpcs.clkbufd3.impl1 analog/buflogic.conv.smpcs.CLKBUFD2
+ AVDD VSS analog/buflogic.conv.smpcs.clkbufd3.Z1 sg13g2f_DEL4
Xanalog/buflogic.conv.smpcs.clkbufd3.impl2 analog/buflogic.conv.smpcs.clkbufd3.Z1
+ AVDD VSS analog/buflogic.conv.smpcs.CLKBUFD3 sg13g2f_BUFFD4
Xanalog/buflogic.conv.smpcs.cpreand.impl analog/buflogic.conv.smpcs.CHOLDB1
+ analog/buflogic.conv.smpcs.CLKBUFD3 AVDD VSS analog/buflogic.PRE
+ sg13g2f_AN2D4
Xanalog/buflogic.conv.smpcs.invsmp.impl SAMPLE AVDD VSS analog/buflogic.HOLD
+ sg13g2f_INVD8
Xanalog/buflogic.lnbuf_ccmp.del4.impl1 analog/buflogic.CMP
+ AVDD VSS analog/buflogic.lnbuf_ccmp.del4.Z1 sg13g2f_DEL4
Xanalog/buflogic.lnbuf_ccmp.del4.impl2 analog/buflogic.lnbuf_ccmp.del4.Z1
+ AVDD VSS analog/buflogic.lnbuf_ccmp.ID sg13g2f_BUFFD4
Xanalog/buflogic.lnbuf_ccmp.deland.impl analog/buflogic.CMP
+ analog/buflogic.lnbuf_ccmp.ID AVDD VSS analog/buflogic.lnbuf_ccmp.IP
+ sg13g2f_AN2D4
Xanalog/buflogic.lnbuf_ccmp.delbuf16.impl analog/buflogic.lnbuf_ccmp.IP
+ AVDD VSS analog/CCMP sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_ccmp.ln1.impl analog/buflogic.CMP AVDD
+ VSS analog/buflogic.lnbuf_ccmp.IL sg13g2f_INVD6
Xanalog/buflogic.lnbuf_ccmp.ln2.impl analog/buflogic.lnbuf_ccmp.IL
+ AVDD VSS analog/buflogic.CMP sg13g2f_INVD6
Xanalog/buflogic.lnbuf_ccmp.lnbbuf16.impl analog/buflogic.lnbuf_ccmp.ILBUF
+ AVDD VSS analog/CCMPB sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_ccmp.lnbbuf4.impl analog/buflogic.lnbuf_ccmp.IL
+ AVDD VSS analog/buflogic.lnbuf_ccmp.ILBUF sg13g2f_BUFFD4
Xanalog/buflogic.lnbuf_chold.ibuf16.impl analog/buflogic.HOLD
+ AVDD VSS analog/buflogic.lnbuf_chold.N3 sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_chold.ln1.impl analog/buflogic.lnbuf_chold.N3
+ AVDD VSS analog/buflogic.lnbuf_chold.N2 sg13g2f_INVD8
Xanalog/buflogic.lnbuf_chold.ln2.impl analog/buflogic.lnbuf_chold.N2
+ AVDD VSS analog/buflogic.lnbuf_chold.N3 sg13g2f_INVD8
Xanalog/buflogic.lnbuf_chold.zbuf16_1.impl analog/buflogic.lnbuf_chold.N1
+ AVDD VSS analog/CHOLD sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_chold.zbuf16_2.impl analog/buflogic.lnbuf_chold.N1
+ AVDD VSS analog/CHOLD sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_chold.zbuf8.impl analog/buflogic.lnbuf_chold.N3
+ AVDD VSS analog/buflogic.lnbuf_chold.N1 sg13g2f_BUFFD8
Xanalog/buflogic.lnbuf_chold.znbuf16_1.impl analog/buflogic.lnbuf_chold.N2
+ AVDD VSS analog/CHOLDB sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_chold.znbuf16_2.impl analog/buflogic.lnbuf_chold.N2
+ AVDD VSS analog/CHOLDB sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_cpre.ibuf16.impl analog/buflogic.PRE
+ AVDD VSS analog/buflogic.lnbuf_cpre.N3 sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_cpre.ln1.impl analog/buflogic.lnbuf_cpre.N3
+ AVDD VSS analog/buflogic.lnbuf_cpre.N2 sg13g2f_INVD8
Xanalog/buflogic.lnbuf_cpre.ln2.impl analog/buflogic.lnbuf_cpre.N2
+ AVDD VSS analog/buflogic.lnbuf_cpre.N3 sg13g2f_INVD8
Xanalog/buflogic.lnbuf_cpre.zbuf16_1.impl analog/buflogic.lnbuf_cpre.N1
+ AVDD VSS analog/CPRE sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_cpre.zbuf16_2.impl analog/buflogic.lnbuf_cpre.N1
+ AVDD VSS analog/CPRE sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_cpre.zbuf8.impl analog/buflogic.lnbuf_cpre.N3
+ AVDD VSS analog/buflogic.lnbuf_cpre.N1 sg13g2f_BUFFD8
Xanalog/buflogic.lnbuf_cpre.znbuf16_1.impl analog/buflogic.lnbuf_cpre.N2
+ AVDD VSS analog/CPREB sg13g2f_BUFFD16
Xanalog/buflogic.lnbuf_cpre.znbuf16_2.impl analog/buflogic.lnbuf_cpre.N2
+ AVDD VSS analog/CPREB sg13g2f_BUFFD16
Xanalog/cmp.buf_n0.impl analog/cmp.OUTNp AVDD VSS analog/cmp.OUTNpb
+ sg13g2f_BUFFD0
Xanalog/cmp.buf_n1.impl analog/cmp.OUTNpb AVDD VSS analog/cmp.OUTN
+ sg13g2f_BUFFD2
Xanalog/cmp.buf_p0.impl analog/cmp.OUTPp AVDD VSS analog/cmp.OUTPpb
+ sg13g2f_BUFFD0
Xanalog/cmp.buf_p1.impl analog/cmp.OUTPpb AVDD VSS CMPO sg13g2f_BUFFD2
Xanalog/cmp.n2p.impl analog/cmp.OUTNp analog/CCMP AVDD VSS
+ analog/cmp.OUTPp sg13g2f_ND2D2
Xanalog/cmp.p2n.impl analog/cmp.OUTPp analog/CCMP AVDD VSS
+ analog/cmp.OUTNp sg13g2f_ND2D2
Xanalog/cmp.vn_cmp.impl_0 analog/CCMPB analog/VOUTL analog/CCMP
+ analog/cmp.OUTNp AVDD VSS analog/cmp.OUTPp sg13g2f_OAI211D4
Xanalog/cmp.vn_cmp.impl_1 analog/CCMPB analog/VOUTL analog/CCMP
+ analog/cmp.OUTNp AVDD VSS analog/cmp.OUTPp sg13g2f_OAI211D4
Xanalog/cmp.vn_cmp.impl_2 analog/CCMPB analog/VOUTL analog/CCMP
+ analog/cmp.OUTNp AVDD VSS analog/cmp.OUTPp sg13g2f_OAI211D4
Xanalog/cmp.vn_cmp.impl_3 analog/CCMPB analog/VOUTL analog/CCMP
+ analog/cmp.OUTNp AVDD VSS analog/cmp.OUTPp sg13g2f_OAI211D4
Xanalog/cmp.vp_cmp.impl_0 analog/CCMPB analog/VOUTH analog/CCMP
+ analog/cmp.OUTPp AVDD VSS analog/cmp.OUTNp sg13g2f_OAI211D4
Xanalog/cmp.vp_cmp.impl_1 analog/CCMPB analog/VOUTH analog/CCMP
+ analog/cmp.OUTPp AVDD VSS analog/cmp.OUTNp sg13g2f_OAI211D4
Xanalog/cmp.vp_cmp.impl_2 analog/CCMPB analog/VOUTH analog/CCMP
+ analog/cmp.OUTPp AVDD VSS analog/cmp.OUTNp sg13g2f_OAI211D4
Xanalog/cmp.vp_cmp.impl_3 analog/CCMPB analog/VOUTH analog/CCMP
+ analog/cmp.OUTPp AVDD VSS analog/cmp.OUTNp sg13g2f_OAI211D4
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[0\].dummy.VSH
+ analog/dummy_h.dummy\[0\].dummy.VOUTH analog/dummy_h.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[0\].dummy.VOUTH
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[0\].dummy.VOUTH
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[0\].dummy.VSH
+ analog/dummy_h.dummy\[0\].dummy.VOUTH analog/dummy_h.dummy\[0\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[0\].dummy.VSH
+ analog/dummy_h.dummy\[0\].dummy.VOUTL analog/dummy_h.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[0\].dummy.VOUTL
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[0\].dummy.VOUTL
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[0\].dummy.VSH
+ analog/dummy_h.dummy\[0\].dummy.VOUTL analog/dummy_h.dummy\[0\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.FL
+ analog/dummy_h.dummy\[0\].dummy.FL analog/dummy_h.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.FL
+ analog/dummy_h.dummy\[0\].dummy.FL analog/dummy_h.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.FL
+ analog/dummy_h.dummy\[0\].dummy.FL analog/dummy_h.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.FL
+ analog/dummy_h.dummy\[0\].dummy.FL analog/dummy_h.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.FL
+ analog/dummy_h.dummy\[0\].dummy.FL analog/dummy_h.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.FL
+ analog/dummy_h.dummy\[0\].dummy.FL analog/dummy_h.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[0\].dummy.VREF
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[0\].dummy.VSH
+ analog/dummy_h.dummy\[0\].dummy.VREF analog/dummy_h.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[0\].dummy.VSH
+ analog/dummy_h.dummy\[0\].dummy.VREF analog/dummy_h.dummy\[0\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[0\].dummy.VREF
+ analog/dummy_h.dummy\[0\].dummy.VSH analog/dummy_h.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[10\].dummy.VSH
+ analog/dummy_h.dummy\[10\].dummy.VOUTH analog/dummy_h.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[10\].dummy.VOUTH
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[10\].dummy.VOUTH
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[10\].dummy.VSH
+ analog/dummy_h.dummy\[10\].dummy.VOUTH analog/dummy_h.dummy\[10\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[10\].dummy.VSH
+ analog/dummy_h.dummy\[10\].dummy.VOUTL analog/dummy_h.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[10\].dummy.VOUTL
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[10\].dummy.VOUTL
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[10\].dummy.VSH
+ analog/dummy_h.dummy\[10\].dummy.VOUTL analog/dummy_h.dummy\[10\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.FL
+ analog/dummy_h.dummy\[10\].dummy.FL analog/dummy_h.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.FL
+ analog/dummy_h.dummy\[10\].dummy.FL analog/dummy_h.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.FL
+ analog/dummy_h.dummy\[10\].dummy.FL analog/dummy_h.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.FL
+ analog/dummy_h.dummy\[10\].dummy.FL analog/dummy_h.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.FL
+ analog/dummy_h.dummy\[10\].dummy.FL analog/dummy_h.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.FL
+ analog/dummy_h.dummy\[10\].dummy.FL analog/dummy_h.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[10\].dummy.VREF
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[10\].dummy.VSH
+ analog/dummy_h.dummy\[10\].dummy.VREF analog/dummy_h.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[10\].dummy.VSH
+ analog/dummy_h.dummy\[10\].dummy.VREF analog/dummy_h.dummy\[10\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[10\].dummy.VREF
+ analog/dummy_h.dummy\[10\].dummy.VSH analog/dummy_h.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[11\].dummy.VSH
+ analog/dummy_h.dummy\[11\].dummy.VOUTH analog/dummy_h.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[11\].dummy.VOUTH
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[11\].dummy.VOUTH
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[11\].dummy.VSH
+ analog/dummy_h.dummy\[11\].dummy.VOUTH analog/dummy_h.dummy\[11\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[11\].dummy.VSH
+ analog/dummy_h.dummy\[11\].dummy.VOUTL analog/dummy_h.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[11\].dummy.VOUTL
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[11\].dummy.VOUTL
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[11\].dummy.VSH
+ analog/dummy_h.dummy\[11\].dummy.VOUTL analog/dummy_h.dummy\[11\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.FL
+ analog/dummy_h.dummy\[11\].dummy.FL analog/dummy_h.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.FL
+ analog/dummy_h.dummy\[11\].dummy.FL analog/dummy_h.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.FL
+ analog/dummy_h.dummy\[11\].dummy.FL analog/dummy_h.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.FL
+ analog/dummy_h.dummy\[11\].dummy.FL analog/dummy_h.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.FL
+ analog/dummy_h.dummy\[11\].dummy.FL analog/dummy_h.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.FL
+ analog/dummy_h.dummy\[11\].dummy.FL analog/dummy_h.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[11\].dummy.VREF
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[11\].dummy.VSH
+ analog/dummy_h.dummy\[11\].dummy.VREF analog/dummy_h.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[11\].dummy.VSH
+ analog/dummy_h.dummy\[11\].dummy.VREF analog/dummy_h.dummy\[11\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[11\].dummy.VREF
+ analog/dummy_h.dummy\[11\].dummy.VSH analog/dummy_h.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[12\].dummy.VSH
+ analog/dummy_h.dummy\[12\].dummy.VOUTH analog/dummy_h.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[12\].dummy.VOUTH
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[12\].dummy.VOUTH
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[12\].dummy.VSH
+ analog/dummy_h.dummy\[12\].dummy.VOUTH analog/dummy_h.dummy\[12\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[12\].dummy.VSH
+ analog/dummy_h.dummy\[12\].dummy.VOUTL analog/dummy_h.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[12\].dummy.VOUTL
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[12\].dummy.VOUTL
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[12\].dummy.VSH
+ analog/dummy_h.dummy\[12\].dummy.VOUTL analog/dummy_h.dummy\[12\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.FL
+ analog/dummy_h.dummy\[12\].dummy.FL analog/dummy_h.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.FL
+ analog/dummy_h.dummy\[12\].dummy.FL analog/dummy_h.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.FL
+ analog/dummy_h.dummy\[12\].dummy.FL analog/dummy_h.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.FL
+ analog/dummy_h.dummy\[12\].dummy.FL analog/dummy_h.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.FL
+ analog/dummy_h.dummy\[12\].dummy.FL analog/dummy_h.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.FL
+ analog/dummy_h.dummy\[12\].dummy.FL analog/dummy_h.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[12\].dummy.VREF
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[12\].dummy.VSH
+ analog/dummy_h.dummy\[12\].dummy.VREF analog/dummy_h.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[12\].dummy.VSH
+ analog/dummy_h.dummy\[12\].dummy.VREF analog/dummy_h.dummy\[12\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[12\].dummy.VREF
+ analog/dummy_h.dummy\[12\].dummy.VSH analog/dummy_h.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[13\].dummy.VSH
+ analog/dummy_h.dummy\[13\].dummy.VOUTH analog/dummy_h.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[13\].dummy.VOUTH
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[13\].dummy.VOUTH
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[13\].dummy.VSH
+ analog/dummy_h.dummy\[13\].dummy.VOUTH analog/dummy_h.dummy\[13\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[13\].dummy.VSH
+ analog/dummy_h.dummy\[13\].dummy.VOUTL analog/dummy_h.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[13\].dummy.VOUTL
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[13\].dummy.VOUTL
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[13\].dummy.VSH
+ analog/dummy_h.dummy\[13\].dummy.VOUTL analog/dummy_h.dummy\[13\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.FL
+ analog/dummy_h.dummy\[13\].dummy.FL analog/dummy_h.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.FL
+ analog/dummy_h.dummy\[13\].dummy.FL analog/dummy_h.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.FL
+ analog/dummy_h.dummy\[13\].dummy.FL analog/dummy_h.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.FL
+ analog/dummy_h.dummy\[13\].dummy.FL analog/dummy_h.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.FL
+ analog/dummy_h.dummy\[13\].dummy.FL analog/dummy_h.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.FL
+ analog/dummy_h.dummy\[13\].dummy.FL analog/dummy_h.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[13\].dummy.VREF
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[13\].dummy.VSH
+ analog/dummy_h.dummy\[13\].dummy.VREF analog/dummy_h.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[13\].dummy.VSH
+ analog/dummy_h.dummy\[13\].dummy.VREF analog/dummy_h.dummy\[13\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[13\].dummy.VREF
+ analog/dummy_h.dummy\[13\].dummy.VSH analog/dummy_h.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[14\].dummy.VSH
+ analog/dummy_h.dummy\[14\].dummy.VOUTH analog/dummy_h.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[14\].dummy.VOUTH
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[14\].dummy.VOUTH
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[14\].dummy.VSH
+ analog/dummy_h.dummy\[14\].dummy.VOUTH analog/dummy_h.dummy\[14\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[14\].dummy.VSH
+ analog/dummy_h.dummy\[14\].dummy.VOUTL analog/dummy_h.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[14\].dummy.VOUTL
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[14\].dummy.VOUTL
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[14\].dummy.VSH
+ analog/dummy_h.dummy\[14\].dummy.VOUTL analog/dummy_h.dummy\[14\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.FL
+ analog/dummy_h.dummy\[14\].dummy.FL analog/dummy_h.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.FL
+ analog/dummy_h.dummy\[14\].dummy.FL analog/dummy_h.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.FL
+ analog/dummy_h.dummy\[14\].dummy.FL analog/dummy_h.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.FL
+ analog/dummy_h.dummy\[14\].dummy.FL analog/dummy_h.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.FL
+ analog/dummy_h.dummy\[14\].dummy.FL analog/dummy_h.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.FL
+ analog/dummy_h.dummy\[14\].dummy.FL analog/dummy_h.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[14\].dummy.VREF
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[14\].dummy.VSH
+ analog/dummy_h.dummy\[14\].dummy.VREF analog/dummy_h.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[14\].dummy.VSH
+ analog/dummy_h.dummy\[14\].dummy.VREF analog/dummy_h.dummy\[14\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[14\].dummy.VREF
+ analog/dummy_h.dummy\[14\].dummy.VSH analog/dummy_h.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[15\].dummy.VSH
+ analog/dummy_h.dummy\[15\].dummy.VOUTH analog/dummy_h.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[15\].dummy.VOUTH
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[15\].dummy.VOUTH
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[15\].dummy.VSH
+ analog/dummy_h.dummy\[15\].dummy.VOUTH analog/dummy_h.dummy\[15\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[15\].dummy.VSH
+ analog/dummy_h.dummy\[15\].dummy.VOUTL analog/dummy_h.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[15\].dummy.VOUTL
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[15\].dummy.VOUTL
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[15\].dummy.VSH
+ analog/dummy_h.dummy\[15\].dummy.VOUTL analog/dummy_h.dummy\[15\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.FL
+ analog/dummy_h.dummy\[15\].dummy.FL analog/dummy_h.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.FL
+ analog/dummy_h.dummy\[15\].dummy.FL analog/dummy_h.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.FL
+ analog/dummy_h.dummy\[15\].dummy.FL analog/dummy_h.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.FL
+ analog/dummy_h.dummy\[15\].dummy.FL analog/dummy_h.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.FL
+ analog/dummy_h.dummy\[15\].dummy.FL analog/dummy_h.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.FL
+ analog/dummy_h.dummy\[15\].dummy.FL analog/dummy_h.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[15\].dummy.VREF
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[15\].dummy.VSH
+ analog/dummy_h.dummy\[15\].dummy.VREF analog/dummy_h.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[15\].dummy.VSH
+ analog/dummy_h.dummy\[15\].dummy.VREF analog/dummy_h.dummy\[15\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[15\].dummy.VREF
+ analog/dummy_h.dummy\[15\].dummy.VSH analog/dummy_h.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[16\].dummy.VSH
+ analog/dummy_h.dummy\[16\].dummy.VOUTH analog/dummy_h.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[16\].dummy.VOUTH
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[16\].dummy.VOUTH
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[16\].dummy.VSH
+ analog/dummy_h.dummy\[16\].dummy.VOUTH analog/dummy_h.dummy\[16\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[16\].dummy.VSH
+ analog/dummy_h.dummy\[16\].dummy.VOUTL analog/dummy_h.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[16\].dummy.VOUTL
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[16\].dummy.VOUTL
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[16\].dummy.VSH
+ analog/dummy_h.dummy\[16\].dummy.VOUTL analog/dummy_h.dummy\[16\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.FL
+ analog/dummy_h.dummy\[16\].dummy.FL analog/dummy_h.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.FL
+ analog/dummy_h.dummy\[16\].dummy.FL analog/dummy_h.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.FL
+ analog/dummy_h.dummy\[16\].dummy.FL analog/dummy_h.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.FL
+ analog/dummy_h.dummy\[16\].dummy.FL analog/dummy_h.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.FL
+ analog/dummy_h.dummy\[16\].dummy.FL analog/dummy_h.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.FL
+ analog/dummy_h.dummy\[16\].dummy.FL analog/dummy_h.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[16\].dummy.VREF
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[16\].dummy.VSH
+ analog/dummy_h.dummy\[16\].dummy.VREF analog/dummy_h.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[16\].dummy.VSH
+ analog/dummy_h.dummy\[16\].dummy.VREF analog/dummy_h.dummy\[16\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[16\].dummy.VREF
+ analog/dummy_h.dummy\[16\].dummy.VSH analog/dummy_h.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[17\].dummy.VSH
+ analog/dummy_h.dummy\[17\].dummy.VOUTH analog/dummy_h.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[17\].dummy.VOUTH
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[17\].dummy.VOUTH
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[17\].dummy.VSH
+ analog/dummy_h.dummy\[17\].dummy.VOUTH analog/dummy_h.dummy\[17\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[17\].dummy.VSH
+ analog/dummy_h.dummy\[17\].dummy.VOUTL analog/dummy_h.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[17\].dummy.VOUTL
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[17\].dummy.VOUTL
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[17\].dummy.VSH
+ analog/dummy_h.dummy\[17\].dummy.VOUTL analog/dummy_h.dummy\[17\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.FL
+ analog/dummy_h.dummy\[17\].dummy.FL analog/dummy_h.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.FL
+ analog/dummy_h.dummy\[17\].dummy.FL analog/dummy_h.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.FL
+ analog/dummy_h.dummy\[17\].dummy.FL analog/dummy_h.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.FL
+ analog/dummy_h.dummy\[17\].dummy.FL analog/dummy_h.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.FL
+ analog/dummy_h.dummy\[17\].dummy.FL analog/dummy_h.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.FL
+ analog/dummy_h.dummy\[17\].dummy.FL analog/dummy_h.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[17\].dummy.VREF
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[17\].dummy.VSH
+ analog/dummy_h.dummy\[17\].dummy.VREF analog/dummy_h.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[17\].dummy.VSH
+ analog/dummy_h.dummy\[17\].dummy.VREF analog/dummy_h.dummy\[17\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[17\].dummy.VREF
+ analog/dummy_h.dummy\[17\].dummy.VSH analog/dummy_h.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[18\].dummy.VSH
+ analog/dummy_h.dummy\[18\].dummy.VOUTH analog/dummy_h.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[18\].dummy.VOUTH
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[18\].dummy.VOUTH
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[18\].dummy.VSH
+ analog/dummy_h.dummy\[18\].dummy.VOUTH analog/dummy_h.dummy\[18\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[18\].dummy.VSH
+ analog/dummy_h.dummy\[18\].dummy.VOUTL analog/dummy_h.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[18\].dummy.VOUTL
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[18\].dummy.VOUTL
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[18\].dummy.VSH
+ analog/dummy_h.dummy\[18\].dummy.VOUTL analog/dummy_h.dummy\[18\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.FL
+ analog/dummy_h.dummy\[18\].dummy.FL analog/dummy_h.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.FL
+ analog/dummy_h.dummy\[18\].dummy.FL analog/dummy_h.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.FL
+ analog/dummy_h.dummy\[18\].dummy.FL analog/dummy_h.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.FL
+ analog/dummy_h.dummy\[18\].dummy.FL analog/dummy_h.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.FL
+ analog/dummy_h.dummy\[18\].dummy.FL analog/dummy_h.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.FL
+ analog/dummy_h.dummy\[18\].dummy.FL analog/dummy_h.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[18\].dummy.VREF
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[18\].dummy.VSH
+ analog/dummy_h.dummy\[18\].dummy.VREF analog/dummy_h.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[18\].dummy.VSH
+ analog/dummy_h.dummy\[18\].dummy.VREF analog/dummy_h.dummy\[18\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[18\].dummy.VREF
+ analog/dummy_h.dummy\[18\].dummy.VSH analog/dummy_h.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[19\].dummy.VSH
+ analog/dummy_h.dummy\[19\].dummy.VOUTH analog/dummy_h.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[19\].dummy.VOUTH
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[19\].dummy.VOUTH
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[19\].dummy.VSH
+ analog/dummy_h.dummy\[19\].dummy.VOUTH analog/dummy_h.dummy\[19\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[19\].dummy.VSH
+ analog/dummy_h.dummy\[19\].dummy.VOUTL analog/dummy_h.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[19\].dummy.VOUTL
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[19\].dummy.VOUTL
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[19\].dummy.VSH
+ analog/dummy_h.dummy\[19\].dummy.VOUTL analog/dummy_h.dummy\[19\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.FL
+ analog/dummy_h.dummy\[19\].dummy.FL analog/dummy_h.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.FL
+ analog/dummy_h.dummy\[19\].dummy.FL analog/dummy_h.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.FL
+ analog/dummy_h.dummy\[19\].dummy.FL analog/dummy_h.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.FL
+ analog/dummy_h.dummy\[19\].dummy.FL analog/dummy_h.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.FL
+ analog/dummy_h.dummy\[19\].dummy.FL analog/dummy_h.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.FL
+ analog/dummy_h.dummy\[19\].dummy.FL analog/dummy_h.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[19\].dummy.VREF
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[19\].dummy.VSH
+ analog/dummy_h.dummy\[19\].dummy.VREF analog/dummy_h.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[19\].dummy.VSH
+ analog/dummy_h.dummy\[19\].dummy.VREF analog/dummy_h.dummy\[19\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[19\].dummy.VREF
+ analog/dummy_h.dummy\[19\].dummy.VSH analog/dummy_h.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[1\].dummy.VSH
+ analog/dummy_h.dummy\[1\].dummy.VOUTH analog/dummy_h.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[1\].dummy.VOUTH
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[1\].dummy.VOUTH
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[1\].dummy.VSH
+ analog/dummy_h.dummy\[1\].dummy.VOUTH analog/dummy_h.dummy\[1\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[1\].dummy.VSH
+ analog/dummy_h.dummy\[1\].dummy.VOUTL analog/dummy_h.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[1\].dummy.VOUTL
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[1\].dummy.VOUTL
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[1\].dummy.VSH
+ analog/dummy_h.dummy\[1\].dummy.VOUTL analog/dummy_h.dummy\[1\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.FL
+ analog/dummy_h.dummy\[1\].dummy.FL analog/dummy_h.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.FL
+ analog/dummy_h.dummy\[1\].dummy.FL analog/dummy_h.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.FL
+ analog/dummy_h.dummy\[1\].dummy.FL analog/dummy_h.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.FL
+ analog/dummy_h.dummy\[1\].dummy.FL analog/dummy_h.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.FL
+ analog/dummy_h.dummy\[1\].dummy.FL analog/dummy_h.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.FL
+ analog/dummy_h.dummy\[1\].dummy.FL analog/dummy_h.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[1\].dummy.VREF
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[1\].dummy.VSH
+ analog/dummy_h.dummy\[1\].dummy.VREF analog/dummy_h.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[1\].dummy.VSH
+ analog/dummy_h.dummy\[1\].dummy.VREF analog/dummy_h.dummy\[1\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[1\].dummy.VREF
+ analog/dummy_h.dummy\[1\].dummy.VSH analog/dummy_h.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[20\].dummy.VSH
+ analog/dummy_h.dummy\[20\].dummy.VOUTH analog/dummy_h.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[20\].dummy.VOUTH
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[20\].dummy.VOUTH
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[20\].dummy.VSH
+ analog/dummy_h.dummy\[20\].dummy.VOUTH analog/dummy_h.dummy\[20\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[20\].dummy.VSH
+ analog/dummy_h.dummy\[20\].dummy.VOUTL analog/dummy_h.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[20\].dummy.VOUTL
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[20\].dummy.VOUTL
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[20\].dummy.VSH
+ analog/dummy_h.dummy\[20\].dummy.VOUTL analog/dummy_h.dummy\[20\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.FL
+ analog/dummy_h.dummy\[20\].dummy.FL analog/dummy_h.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.FL
+ analog/dummy_h.dummy\[20\].dummy.FL analog/dummy_h.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.FL
+ analog/dummy_h.dummy\[20\].dummy.FL analog/dummy_h.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.FL
+ analog/dummy_h.dummy\[20\].dummy.FL analog/dummy_h.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.FL
+ analog/dummy_h.dummy\[20\].dummy.FL analog/dummy_h.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.FL
+ analog/dummy_h.dummy\[20\].dummy.FL analog/dummy_h.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[20\].dummy.VREF
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[20\].dummy.VSH
+ analog/dummy_h.dummy\[20\].dummy.VREF analog/dummy_h.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[20\].dummy.VSH
+ analog/dummy_h.dummy\[20\].dummy.VREF analog/dummy_h.dummy\[20\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[20\].dummy.VREF
+ analog/dummy_h.dummy\[20\].dummy.VSH analog/dummy_h.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[21\].dummy.VSH
+ analog/dummy_h.dummy\[21\].dummy.VOUTH analog/dummy_h.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[21\].dummy.VOUTH
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[21\].dummy.VOUTH
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[21\].dummy.VSH
+ analog/dummy_h.dummy\[21\].dummy.VOUTH analog/dummy_h.dummy\[21\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[21\].dummy.VSH
+ analog/dummy_h.dummy\[21\].dummy.VOUTL analog/dummy_h.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[21\].dummy.VOUTL
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[21\].dummy.VOUTL
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[21\].dummy.VSH
+ analog/dummy_h.dummy\[21\].dummy.VOUTL analog/dummy_h.dummy\[21\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.FL
+ analog/dummy_h.dummy\[21\].dummy.FL analog/dummy_h.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.FL
+ analog/dummy_h.dummy\[21\].dummy.FL analog/dummy_h.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.FL
+ analog/dummy_h.dummy\[21\].dummy.FL analog/dummy_h.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.FL
+ analog/dummy_h.dummy\[21\].dummy.FL analog/dummy_h.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.FL
+ analog/dummy_h.dummy\[21\].dummy.FL analog/dummy_h.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.FL
+ analog/dummy_h.dummy\[21\].dummy.FL analog/dummy_h.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[21\].dummy.VREF
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[21\].dummy.VSH
+ analog/dummy_h.dummy\[21\].dummy.VREF analog/dummy_h.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[21\].dummy.VSH
+ analog/dummy_h.dummy\[21\].dummy.VREF analog/dummy_h.dummy\[21\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[21\].dummy.VREF
+ analog/dummy_h.dummy\[21\].dummy.VSH analog/dummy_h.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[22\].dummy.VSH
+ analog/dummy_h.dummy\[22\].dummy.VOUTH analog/dummy_h.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[22\].dummy.VOUTH
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[22\].dummy.VOUTH
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[22\].dummy.VSH
+ analog/dummy_h.dummy\[22\].dummy.VOUTH analog/dummy_h.dummy\[22\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[22\].dummy.VSH
+ analog/dummy_h.dummy\[22\].dummy.VOUTL analog/dummy_h.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[22\].dummy.VOUTL
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[22\].dummy.VOUTL
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[22\].dummy.VSH
+ analog/dummy_h.dummy\[22\].dummy.VOUTL analog/dummy_h.dummy\[22\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.FL
+ analog/dummy_h.dummy\[22\].dummy.FL analog/dummy_h.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.FL
+ analog/dummy_h.dummy\[22\].dummy.FL analog/dummy_h.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.FL
+ analog/dummy_h.dummy\[22\].dummy.FL analog/dummy_h.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.FL
+ analog/dummy_h.dummy\[22\].dummy.FL analog/dummy_h.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.FL
+ analog/dummy_h.dummy\[22\].dummy.FL analog/dummy_h.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.FL
+ analog/dummy_h.dummy\[22\].dummy.FL analog/dummy_h.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[22\].dummy.VREF
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[22\].dummy.VSH
+ analog/dummy_h.dummy\[22\].dummy.VREF analog/dummy_h.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[22\].dummy.VSH
+ analog/dummy_h.dummy\[22\].dummy.VREF analog/dummy_h.dummy\[22\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[22\].dummy.VREF
+ analog/dummy_h.dummy\[22\].dummy.VSH analog/dummy_h.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[23\].dummy.VSH
+ analog/dummy_h.dummy\[23\].dummy.VOUTH analog/dummy_h.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[23\].dummy.VOUTH
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[23\].dummy.VOUTH
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[23\].dummy.VSH
+ analog/dummy_h.dummy\[23\].dummy.VOUTH analog/dummy_h.dummy\[23\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[23\].dummy.VSH
+ analog/dummy_h.dummy\[23\].dummy.VOUTL analog/dummy_h.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[23\].dummy.VOUTL
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[23\].dummy.VOUTL
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[23\].dummy.VSH
+ analog/dummy_h.dummy\[23\].dummy.VOUTL analog/dummy_h.dummy\[23\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.FL
+ analog/dummy_h.dummy\[23\].dummy.FL analog/dummy_h.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.FL
+ analog/dummy_h.dummy\[23\].dummy.FL analog/dummy_h.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.FL
+ analog/dummy_h.dummy\[23\].dummy.FL analog/dummy_h.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.FL
+ analog/dummy_h.dummy\[23\].dummy.FL analog/dummy_h.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.FL
+ analog/dummy_h.dummy\[23\].dummy.FL analog/dummy_h.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.FL
+ analog/dummy_h.dummy\[23\].dummy.FL analog/dummy_h.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[23\].dummy.VREF
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[23\].dummy.VSH
+ analog/dummy_h.dummy\[23\].dummy.VREF analog/dummy_h.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[23\].dummy.VSH
+ analog/dummy_h.dummy\[23\].dummy.VREF analog/dummy_h.dummy\[23\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[23\].dummy.VREF
+ analog/dummy_h.dummy\[23\].dummy.VSH analog/dummy_h.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[24\].dummy.VSH
+ analog/dummy_h.dummy\[24\].dummy.VOUTH analog/dummy_h.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[24\].dummy.VOUTH
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[24\].dummy.VOUTH
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[24\].dummy.VSH
+ analog/dummy_h.dummy\[24\].dummy.VOUTH analog/dummy_h.dummy\[24\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[24\].dummy.VSH
+ analog/dummy_h.dummy\[24\].dummy.VOUTL analog/dummy_h.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[24\].dummy.VOUTL
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[24\].dummy.VOUTL
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[24\].dummy.VSH
+ analog/dummy_h.dummy\[24\].dummy.VOUTL analog/dummy_h.dummy\[24\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.FL
+ analog/dummy_h.dummy\[24\].dummy.FL analog/dummy_h.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.FL
+ analog/dummy_h.dummy\[24\].dummy.FL analog/dummy_h.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.FL
+ analog/dummy_h.dummy\[24\].dummy.FL analog/dummy_h.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.FL
+ analog/dummy_h.dummy\[24\].dummy.FL analog/dummy_h.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.FL
+ analog/dummy_h.dummy\[24\].dummy.FL analog/dummy_h.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.FL
+ analog/dummy_h.dummy\[24\].dummy.FL analog/dummy_h.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[24\].dummy.VREF
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[24\].dummy.VSH
+ analog/dummy_h.dummy\[24\].dummy.VREF analog/dummy_h.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[24\].dummy.VSH
+ analog/dummy_h.dummy\[24\].dummy.VREF analog/dummy_h.dummy\[24\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[24\].dummy.VREF
+ analog/dummy_h.dummy\[24\].dummy.VSH analog/dummy_h.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[25\].dummy.VSH
+ analog/dummy_h.dummy\[25\].dummy.VOUTH analog/dummy_h.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[25\].dummy.VOUTH
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[25\].dummy.VOUTH
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[25\].dummy.VSH
+ analog/dummy_h.dummy\[25\].dummy.VOUTH analog/dummy_h.dummy\[25\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[25\].dummy.VSH
+ analog/dummy_h.dummy\[25\].dummy.VOUTL analog/dummy_h.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[25\].dummy.VOUTL
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[25\].dummy.VOUTL
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[25\].dummy.VSH
+ analog/dummy_h.dummy\[25\].dummy.VOUTL analog/dummy_h.dummy\[25\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.FL
+ analog/dummy_h.dummy\[25\].dummy.FL analog/dummy_h.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.FL
+ analog/dummy_h.dummy\[25\].dummy.FL analog/dummy_h.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.FL
+ analog/dummy_h.dummy\[25\].dummy.FL analog/dummy_h.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.FL
+ analog/dummy_h.dummy\[25\].dummy.FL analog/dummy_h.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.FL
+ analog/dummy_h.dummy\[25\].dummy.FL analog/dummy_h.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.FL
+ analog/dummy_h.dummy\[25\].dummy.FL analog/dummy_h.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[25\].dummy.VREF
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[25\].dummy.VSH
+ analog/dummy_h.dummy\[25\].dummy.VREF analog/dummy_h.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[25\].dummy.VSH
+ analog/dummy_h.dummy\[25\].dummy.VREF analog/dummy_h.dummy\[25\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[25\].dummy.VREF
+ analog/dummy_h.dummy\[25\].dummy.VSH analog/dummy_h.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[26\].dummy.VSH
+ analog/dummy_h.dummy\[26\].dummy.VOUTH analog/dummy_h.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[26\].dummy.VOUTH
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[26\].dummy.VOUTH
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[26\].dummy.VSH
+ analog/dummy_h.dummy\[26\].dummy.VOUTH analog/dummy_h.dummy\[26\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[26\].dummy.VSH
+ analog/dummy_h.dummy\[26\].dummy.VOUTL analog/dummy_h.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[26\].dummy.VOUTL
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[26\].dummy.VOUTL
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[26\].dummy.VSH
+ analog/dummy_h.dummy\[26\].dummy.VOUTL analog/dummy_h.dummy\[26\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.FL
+ analog/dummy_h.dummy\[26\].dummy.FL analog/dummy_h.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.FL
+ analog/dummy_h.dummy\[26\].dummy.FL analog/dummy_h.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.FL
+ analog/dummy_h.dummy\[26\].dummy.FL analog/dummy_h.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.FL
+ analog/dummy_h.dummy\[26\].dummy.FL analog/dummy_h.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.FL
+ analog/dummy_h.dummy\[26\].dummy.FL analog/dummy_h.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.FL
+ analog/dummy_h.dummy\[26\].dummy.FL analog/dummy_h.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[26\].dummy.VREF
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[26\].dummy.VSH
+ analog/dummy_h.dummy\[26\].dummy.VREF analog/dummy_h.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[26\].dummy.VSH
+ analog/dummy_h.dummy\[26\].dummy.VREF analog/dummy_h.dummy\[26\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[26\].dummy.VREF
+ analog/dummy_h.dummy\[26\].dummy.VSH analog/dummy_h.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[27\].dummy.VSH
+ analog/dummy_h.dummy\[27\].dummy.VOUTH analog/dummy_h.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[27\].dummy.VOUTH
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[27\].dummy.VOUTH
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[27\].dummy.VSH
+ analog/dummy_h.dummy\[27\].dummy.VOUTH analog/dummy_h.dummy\[27\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[27\].dummy.VSH
+ analog/dummy_h.dummy\[27\].dummy.VOUTL analog/dummy_h.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[27\].dummy.VOUTL
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[27\].dummy.VOUTL
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[27\].dummy.VSH
+ analog/dummy_h.dummy\[27\].dummy.VOUTL analog/dummy_h.dummy\[27\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.FL
+ analog/dummy_h.dummy\[27\].dummy.FL analog/dummy_h.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.FL
+ analog/dummy_h.dummy\[27\].dummy.FL analog/dummy_h.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.FL
+ analog/dummy_h.dummy\[27\].dummy.FL analog/dummy_h.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.FL
+ analog/dummy_h.dummy\[27\].dummy.FL analog/dummy_h.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.FL
+ analog/dummy_h.dummy\[27\].dummy.FL analog/dummy_h.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.FL
+ analog/dummy_h.dummy\[27\].dummy.FL analog/dummy_h.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[27\].dummy.VREF
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[27\].dummy.VSH
+ analog/dummy_h.dummy\[27\].dummy.VREF analog/dummy_h.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[27\].dummy.VSH
+ analog/dummy_h.dummy\[27\].dummy.VREF analog/dummy_h.dummy\[27\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[27\].dummy.VREF
+ analog/dummy_h.dummy\[27\].dummy.VSH analog/dummy_h.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[2\].dummy.VSH
+ analog/dummy_h.dummy\[2\].dummy.VOUTH analog/dummy_h.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[2\].dummy.VOUTH
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[2\].dummy.VOUTH
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[2\].dummy.VSH
+ analog/dummy_h.dummy\[2\].dummy.VOUTH analog/dummy_h.dummy\[2\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[2\].dummy.VSH
+ analog/dummy_h.dummy\[2\].dummy.VOUTL analog/dummy_h.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[2\].dummy.VOUTL
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[2\].dummy.VOUTL
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[2\].dummy.VSH
+ analog/dummy_h.dummy\[2\].dummy.VOUTL analog/dummy_h.dummy\[2\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.FL
+ analog/dummy_h.dummy\[2\].dummy.FL analog/dummy_h.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.FL
+ analog/dummy_h.dummy\[2\].dummy.FL analog/dummy_h.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.FL
+ analog/dummy_h.dummy\[2\].dummy.FL analog/dummy_h.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.FL
+ analog/dummy_h.dummy\[2\].dummy.FL analog/dummy_h.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.FL
+ analog/dummy_h.dummy\[2\].dummy.FL analog/dummy_h.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.FL
+ analog/dummy_h.dummy\[2\].dummy.FL analog/dummy_h.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[2\].dummy.VREF
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[2\].dummy.VSH
+ analog/dummy_h.dummy\[2\].dummy.VREF analog/dummy_h.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[2\].dummy.VSH
+ analog/dummy_h.dummy\[2\].dummy.VREF analog/dummy_h.dummy\[2\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[2\].dummy.VREF
+ analog/dummy_h.dummy\[2\].dummy.VSH analog/dummy_h.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[3\].dummy.VSH
+ analog/dummy_h.dummy\[3\].dummy.VOUTH analog/dummy_h.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[3\].dummy.VOUTH
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[3\].dummy.VOUTH
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[3\].dummy.VSH
+ analog/dummy_h.dummy\[3\].dummy.VOUTH analog/dummy_h.dummy\[3\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[3\].dummy.VSH
+ analog/dummy_h.dummy\[3\].dummy.VOUTL analog/dummy_h.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[3\].dummy.VOUTL
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[3\].dummy.VOUTL
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[3\].dummy.VSH
+ analog/dummy_h.dummy\[3\].dummy.VOUTL analog/dummy_h.dummy\[3\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.FL
+ analog/dummy_h.dummy\[3\].dummy.FL analog/dummy_h.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.FL
+ analog/dummy_h.dummy\[3\].dummy.FL analog/dummy_h.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.FL
+ analog/dummy_h.dummy\[3\].dummy.FL analog/dummy_h.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.FL
+ analog/dummy_h.dummy\[3\].dummy.FL analog/dummy_h.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.FL
+ analog/dummy_h.dummy\[3\].dummy.FL analog/dummy_h.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.FL
+ analog/dummy_h.dummy\[3\].dummy.FL analog/dummy_h.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[3\].dummy.VREF
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[3\].dummy.VSH
+ analog/dummy_h.dummy\[3\].dummy.VREF analog/dummy_h.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[3\].dummy.VSH
+ analog/dummy_h.dummy\[3\].dummy.VREF analog/dummy_h.dummy\[3\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[3\].dummy.VREF
+ analog/dummy_h.dummy\[3\].dummy.VSH analog/dummy_h.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[4\].dummy.VSH
+ analog/dummy_h.dummy\[4\].dummy.VOUTH analog/dummy_h.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[4\].dummy.VOUTH
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[4\].dummy.VOUTH
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[4\].dummy.VSH
+ analog/dummy_h.dummy\[4\].dummy.VOUTH analog/dummy_h.dummy\[4\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[4\].dummy.VSH
+ analog/dummy_h.dummy\[4\].dummy.VOUTL analog/dummy_h.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[4\].dummy.VOUTL
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[4\].dummy.VOUTL
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[4\].dummy.VSH
+ analog/dummy_h.dummy\[4\].dummy.VOUTL analog/dummy_h.dummy\[4\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.FL
+ analog/dummy_h.dummy\[4\].dummy.FL analog/dummy_h.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.FL
+ analog/dummy_h.dummy\[4\].dummy.FL analog/dummy_h.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.FL
+ analog/dummy_h.dummy\[4\].dummy.FL analog/dummy_h.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.FL
+ analog/dummy_h.dummy\[4\].dummy.FL analog/dummy_h.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.FL
+ analog/dummy_h.dummy\[4\].dummy.FL analog/dummy_h.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.FL
+ analog/dummy_h.dummy\[4\].dummy.FL analog/dummy_h.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[4\].dummy.VREF
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[4\].dummy.VSH
+ analog/dummy_h.dummy\[4\].dummy.VREF analog/dummy_h.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[4\].dummy.VSH
+ analog/dummy_h.dummy\[4\].dummy.VREF analog/dummy_h.dummy\[4\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[4\].dummy.VREF
+ analog/dummy_h.dummy\[4\].dummy.VSH analog/dummy_h.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[5\].dummy.VSH
+ analog/dummy_h.dummy\[5\].dummy.VOUTH analog/dummy_h.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[5\].dummy.VOUTH
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[5\].dummy.VOUTH
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[5\].dummy.VSH
+ analog/dummy_h.dummy\[5\].dummy.VOUTH analog/dummy_h.dummy\[5\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[5\].dummy.VSH
+ analog/dummy_h.dummy\[5\].dummy.VOUTL analog/dummy_h.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[5\].dummy.VOUTL
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[5\].dummy.VOUTL
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[5\].dummy.VSH
+ analog/dummy_h.dummy\[5\].dummy.VOUTL analog/dummy_h.dummy\[5\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.FL
+ analog/dummy_h.dummy\[5\].dummy.FL analog/dummy_h.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.FL
+ analog/dummy_h.dummy\[5\].dummy.FL analog/dummy_h.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.FL
+ analog/dummy_h.dummy\[5\].dummy.FL analog/dummy_h.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.FL
+ analog/dummy_h.dummy\[5\].dummy.FL analog/dummy_h.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.FL
+ analog/dummy_h.dummy\[5\].dummy.FL analog/dummy_h.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.FL
+ analog/dummy_h.dummy\[5\].dummy.FL analog/dummy_h.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[5\].dummy.VREF
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[5\].dummy.VSH
+ analog/dummy_h.dummy\[5\].dummy.VREF analog/dummy_h.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[5\].dummy.VSH
+ analog/dummy_h.dummy\[5\].dummy.VREF analog/dummy_h.dummy\[5\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[5\].dummy.VREF
+ analog/dummy_h.dummy\[5\].dummy.VSH analog/dummy_h.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[6\].dummy.VSH
+ analog/dummy_h.dummy\[6\].dummy.VOUTH analog/dummy_h.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[6\].dummy.VOUTH
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[6\].dummy.VOUTH
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[6\].dummy.VSH
+ analog/dummy_h.dummy\[6\].dummy.VOUTH analog/dummy_h.dummy\[6\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[6\].dummy.VSH
+ analog/dummy_h.dummy\[6\].dummy.VOUTL analog/dummy_h.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[6\].dummy.VOUTL
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[6\].dummy.VOUTL
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[6\].dummy.VSH
+ analog/dummy_h.dummy\[6\].dummy.VOUTL analog/dummy_h.dummy\[6\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.FL
+ analog/dummy_h.dummy\[6\].dummy.FL analog/dummy_h.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.FL
+ analog/dummy_h.dummy\[6\].dummy.FL analog/dummy_h.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.FL
+ analog/dummy_h.dummy\[6\].dummy.FL analog/dummy_h.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.FL
+ analog/dummy_h.dummy\[6\].dummy.FL analog/dummy_h.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.FL
+ analog/dummy_h.dummy\[6\].dummy.FL analog/dummy_h.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.FL
+ analog/dummy_h.dummy\[6\].dummy.FL analog/dummy_h.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[6\].dummy.VREF
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[6\].dummy.VSH
+ analog/dummy_h.dummy\[6\].dummy.VREF analog/dummy_h.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[6\].dummy.VSH
+ analog/dummy_h.dummy\[6\].dummy.VREF analog/dummy_h.dummy\[6\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[6\].dummy.VREF
+ analog/dummy_h.dummy\[6\].dummy.VSH analog/dummy_h.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[7\].dummy.VSH
+ analog/dummy_h.dummy\[7\].dummy.VOUTH analog/dummy_h.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[7\].dummy.VOUTH
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[7\].dummy.VOUTH
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[7\].dummy.VSH
+ analog/dummy_h.dummy\[7\].dummy.VOUTH analog/dummy_h.dummy\[7\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[7\].dummy.VSH
+ analog/dummy_h.dummy\[7\].dummy.VOUTL analog/dummy_h.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[7\].dummy.VOUTL
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[7\].dummy.VOUTL
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[7\].dummy.VSH
+ analog/dummy_h.dummy\[7\].dummy.VOUTL analog/dummy_h.dummy\[7\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.FL
+ analog/dummy_h.dummy\[7\].dummy.FL analog/dummy_h.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.FL
+ analog/dummy_h.dummy\[7\].dummy.FL analog/dummy_h.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.FL
+ analog/dummy_h.dummy\[7\].dummy.FL analog/dummy_h.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.FL
+ analog/dummy_h.dummy\[7\].dummy.FL analog/dummy_h.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.FL
+ analog/dummy_h.dummy\[7\].dummy.FL analog/dummy_h.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.FL
+ analog/dummy_h.dummy\[7\].dummy.FL analog/dummy_h.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[7\].dummy.VREF
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[7\].dummy.VSH
+ analog/dummy_h.dummy\[7\].dummy.VREF analog/dummy_h.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[7\].dummy.VSH
+ analog/dummy_h.dummy\[7\].dummy.VREF analog/dummy_h.dummy\[7\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[7\].dummy.VREF
+ analog/dummy_h.dummy\[7\].dummy.VSH analog/dummy_h.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[8\].dummy.VSH
+ analog/dummy_h.dummy\[8\].dummy.VOUTH analog/dummy_h.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[8\].dummy.VOUTH
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[8\].dummy.VOUTH
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[8\].dummy.VSH
+ analog/dummy_h.dummy\[8\].dummy.VOUTH analog/dummy_h.dummy\[8\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[8\].dummy.VSH
+ analog/dummy_h.dummy\[8\].dummy.VOUTL analog/dummy_h.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[8\].dummy.VOUTL
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[8\].dummy.VOUTL
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[8\].dummy.VSH
+ analog/dummy_h.dummy\[8\].dummy.VOUTL analog/dummy_h.dummy\[8\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.FL
+ analog/dummy_h.dummy\[8\].dummy.FL analog/dummy_h.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.FL
+ analog/dummy_h.dummy\[8\].dummy.FL analog/dummy_h.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.FL
+ analog/dummy_h.dummy\[8\].dummy.FL analog/dummy_h.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.FL
+ analog/dummy_h.dummy\[8\].dummy.FL analog/dummy_h.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.FL
+ analog/dummy_h.dummy\[8\].dummy.FL analog/dummy_h.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.FL
+ analog/dummy_h.dummy\[8\].dummy.FL analog/dummy_h.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[8\].dummy.VREF
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[8\].dummy.VSH
+ analog/dummy_h.dummy\[8\].dummy.VREF analog/dummy_h.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[8\].dummy.VSH
+ analog/dummy_h.dummy\[8\].dummy.VREF analog/dummy_h.dummy\[8\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[8\].dummy.VREF
+ analog/dummy_h.dummy\[8\].dummy.VSH analog/dummy_h.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[9\].dummy.VSH
+ analog/dummy_h.dummy\[9\].dummy.VOUTH analog/dummy_h.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[9\].dummy.VOUTH
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[9\].dummy.VOUTH
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[9\].dummy.VSH
+ analog/dummy_h.dummy\[9\].dummy.VOUTH analog/dummy_h.dummy\[9\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[9\].dummy.VSH
+ analog/dummy_h.dummy\[9\].dummy.VOUTL analog/dummy_h.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[9\].dummy.VOUTL
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[9\].dummy.VOUTL
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[9\].dummy.VSH
+ analog/dummy_h.dummy\[9\].dummy.VOUTL analog/dummy_h.dummy\[9\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.FL
+ analog/dummy_h.dummy\[9\].dummy.FL analog/dummy_h.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.FL
+ analog/dummy_h.dummy\[9\].dummy.FL analog/dummy_h.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.FL
+ analog/dummy_h.dummy\[9\].dummy.FL analog/dummy_h.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.FL
+ analog/dummy_h.dummy\[9\].dummy.FL analog/dummy_h.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.FL
+ analog/dummy_h.dummy\[9\].dummy.FL analog/dummy_h.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.FL
+ analog/dummy_h.dummy\[9\].dummy.FL analog/dummy_h.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[9\].dummy.VREF
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRH analog/dummy_h.dummy\[9\].dummy.VSH
+ analog/dummy_h.dummy\[9\].dummy.VREF analog/dummy_h.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[9\].dummy.VSH
+ analog/dummy_h.dummy\[9\].dummy.VREF analog/dummy_h.dummy\[9\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_h.dummy\[0\].dummy.CRHB analog/dummy_h.dummy\[9\].dummy.VREF
+ analog/dummy_h.dummy\[9\].dummy.VSH analog/dummy_h.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_h.tieh.impl AVDD VSS analog/dummy_h.dummy\[0\].dummy.CRHB
+ sg13g2f_TIEH
Xanalog/dummy_h.tiel.impl AVDD VSS analog/dummy_h.dummy\[0\].dummy.CRH
+ sg13g2f_TIEL
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[0\].dummy.VSH
+ analog/dummy_l.dummy\[0\].dummy.VOUTH analog/dummy_l.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[0\].dummy.VOUTH
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[0\].dummy.VOUTH
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[0\].dummy.VSH
+ analog/dummy_l.dummy\[0\].dummy.VOUTH analog/dummy_l.dummy\[0\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[0\].dummy.VSH
+ analog/dummy_l.dummy\[0\].dummy.VOUTL analog/dummy_l.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[0\].dummy.VOUTL
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[0\].dummy.VOUTL
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[0\].dummy.VSH
+ analog/dummy_l.dummy\[0\].dummy.VOUTL analog/dummy_l.dummy\[0\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.FL
+ analog/dummy_l.dummy\[0\].dummy.FL analog/dummy_l.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.FL
+ analog/dummy_l.dummy\[0\].dummy.FL analog/dummy_l.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.FL
+ analog/dummy_l.dummy\[0\].dummy.FL analog/dummy_l.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.FL
+ analog/dummy_l.dummy\[0\].dummy.FL analog/dummy_l.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.FL
+ analog/dummy_l.dummy\[0\].dummy.FL analog/dummy_l.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.FL
+ analog/dummy_l.dummy\[0\].dummy.FL analog/dummy_l.dummy\[0\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[0\].dummy.VREF
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[0\].dummy.VSH
+ analog/dummy_l.dummy\[0\].dummy.VREF analog/dummy_l.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[0\].dummy.VSH
+ analog/dummy_l.dummy\[0\].dummy.VREF analog/dummy_l.dummy\[0\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[0\].dummy.VREF
+ analog/dummy_l.dummy\[0\].dummy.VSH analog/dummy_l.dummy\[0\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[10\].dummy.VSH
+ analog/dummy_l.dummy\[10\].dummy.VOUTH analog/dummy_l.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[10\].dummy.VOUTH
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[10\].dummy.VOUTH
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[10\].dummy.VSH
+ analog/dummy_l.dummy\[10\].dummy.VOUTH analog/dummy_l.dummy\[10\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[10\].dummy.VSH
+ analog/dummy_l.dummy\[10\].dummy.VOUTL analog/dummy_l.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[10\].dummy.VOUTL
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[10\].dummy.VOUTL
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[10\].dummy.VSH
+ analog/dummy_l.dummy\[10\].dummy.VOUTL analog/dummy_l.dummy\[10\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.FL
+ analog/dummy_l.dummy\[10\].dummy.FL analog/dummy_l.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.FL
+ analog/dummy_l.dummy\[10\].dummy.FL analog/dummy_l.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.FL
+ analog/dummy_l.dummy\[10\].dummy.FL analog/dummy_l.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.FL
+ analog/dummy_l.dummy\[10\].dummy.FL analog/dummy_l.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.FL
+ analog/dummy_l.dummy\[10\].dummy.FL analog/dummy_l.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.FL
+ analog/dummy_l.dummy\[10\].dummy.FL analog/dummy_l.dummy\[10\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[10\].dummy.VREF
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[10\].dummy.VSH
+ analog/dummy_l.dummy\[10\].dummy.VREF analog/dummy_l.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[10\].dummy.VSH
+ analog/dummy_l.dummy\[10\].dummy.VREF analog/dummy_l.dummy\[10\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[10\].dummy.VREF
+ analog/dummy_l.dummy\[10\].dummy.VSH analog/dummy_l.dummy\[10\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[11\].dummy.VSH
+ analog/dummy_l.dummy\[11\].dummy.VOUTH analog/dummy_l.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[11\].dummy.VOUTH
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[11\].dummy.VOUTH
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[11\].dummy.VSH
+ analog/dummy_l.dummy\[11\].dummy.VOUTH analog/dummy_l.dummy\[11\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[11\].dummy.VSH
+ analog/dummy_l.dummy\[11\].dummy.VOUTL analog/dummy_l.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[11\].dummy.VOUTL
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[11\].dummy.VOUTL
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[11\].dummy.VSH
+ analog/dummy_l.dummy\[11\].dummy.VOUTL analog/dummy_l.dummy\[11\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.FL
+ analog/dummy_l.dummy\[11\].dummy.FL analog/dummy_l.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.FL
+ analog/dummy_l.dummy\[11\].dummy.FL analog/dummy_l.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.FL
+ analog/dummy_l.dummy\[11\].dummy.FL analog/dummy_l.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.FL
+ analog/dummy_l.dummy\[11\].dummy.FL analog/dummy_l.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.FL
+ analog/dummy_l.dummy\[11\].dummy.FL analog/dummy_l.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.FL
+ analog/dummy_l.dummy\[11\].dummy.FL analog/dummy_l.dummy\[11\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[11\].dummy.VREF
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[11\].dummy.VSH
+ analog/dummy_l.dummy\[11\].dummy.VREF analog/dummy_l.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[11\].dummy.VSH
+ analog/dummy_l.dummy\[11\].dummy.VREF analog/dummy_l.dummy\[11\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[11\].dummy.VREF
+ analog/dummy_l.dummy\[11\].dummy.VSH analog/dummy_l.dummy\[11\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[12\].dummy.VSH
+ analog/dummy_l.dummy\[12\].dummy.VOUTH analog/dummy_l.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[12\].dummy.VOUTH
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[12\].dummy.VOUTH
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[12\].dummy.VSH
+ analog/dummy_l.dummy\[12\].dummy.VOUTH analog/dummy_l.dummy\[12\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[12\].dummy.VSH
+ analog/dummy_l.dummy\[12\].dummy.VOUTL analog/dummy_l.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[12\].dummy.VOUTL
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[12\].dummy.VOUTL
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[12\].dummy.VSH
+ analog/dummy_l.dummy\[12\].dummy.VOUTL analog/dummy_l.dummy\[12\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.FL
+ analog/dummy_l.dummy\[12\].dummy.FL analog/dummy_l.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.FL
+ analog/dummy_l.dummy\[12\].dummy.FL analog/dummy_l.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.FL
+ analog/dummy_l.dummy\[12\].dummy.FL analog/dummy_l.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.FL
+ analog/dummy_l.dummy\[12\].dummy.FL analog/dummy_l.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.FL
+ analog/dummy_l.dummy\[12\].dummy.FL analog/dummy_l.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.FL
+ analog/dummy_l.dummy\[12\].dummy.FL analog/dummy_l.dummy\[12\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[12\].dummy.VREF
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[12\].dummy.VSH
+ analog/dummy_l.dummy\[12\].dummy.VREF analog/dummy_l.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[12\].dummy.VSH
+ analog/dummy_l.dummy\[12\].dummy.VREF analog/dummy_l.dummy\[12\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[12\].dummy.VREF
+ analog/dummy_l.dummy\[12\].dummy.VSH analog/dummy_l.dummy\[12\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[13\].dummy.VSH
+ analog/dummy_l.dummy\[13\].dummy.VOUTH analog/dummy_l.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[13\].dummy.VOUTH
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[13\].dummy.VOUTH
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[13\].dummy.VSH
+ analog/dummy_l.dummy\[13\].dummy.VOUTH analog/dummy_l.dummy\[13\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[13\].dummy.VSH
+ analog/dummy_l.dummy\[13\].dummy.VOUTL analog/dummy_l.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[13\].dummy.VOUTL
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[13\].dummy.VOUTL
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[13\].dummy.VSH
+ analog/dummy_l.dummy\[13\].dummy.VOUTL analog/dummy_l.dummy\[13\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.FL
+ analog/dummy_l.dummy\[13\].dummy.FL analog/dummy_l.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.FL
+ analog/dummy_l.dummy\[13\].dummy.FL analog/dummy_l.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.FL
+ analog/dummy_l.dummy\[13\].dummy.FL analog/dummy_l.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.FL
+ analog/dummy_l.dummy\[13\].dummy.FL analog/dummy_l.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.FL
+ analog/dummy_l.dummy\[13\].dummy.FL analog/dummy_l.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.FL
+ analog/dummy_l.dummy\[13\].dummy.FL analog/dummy_l.dummy\[13\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[13\].dummy.VREF
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[13\].dummy.VSH
+ analog/dummy_l.dummy\[13\].dummy.VREF analog/dummy_l.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[13\].dummy.VSH
+ analog/dummy_l.dummy\[13\].dummy.VREF analog/dummy_l.dummy\[13\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[13\].dummy.VREF
+ analog/dummy_l.dummy\[13\].dummy.VSH analog/dummy_l.dummy\[13\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[14\].dummy.VSH
+ analog/dummy_l.dummy\[14\].dummy.VOUTH analog/dummy_l.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[14\].dummy.VOUTH
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[14\].dummy.VOUTH
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[14\].dummy.VSH
+ analog/dummy_l.dummy\[14\].dummy.VOUTH analog/dummy_l.dummy\[14\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[14\].dummy.VSH
+ analog/dummy_l.dummy\[14\].dummy.VOUTL analog/dummy_l.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[14\].dummy.VOUTL
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[14\].dummy.VOUTL
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[14\].dummy.VSH
+ analog/dummy_l.dummy\[14\].dummy.VOUTL analog/dummy_l.dummy\[14\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.FL
+ analog/dummy_l.dummy\[14\].dummy.FL analog/dummy_l.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.FL
+ analog/dummy_l.dummy\[14\].dummy.FL analog/dummy_l.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.FL
+ analog/dummy_l.dummy\[14\].dummy.FL analog/dummy_l.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.FL
+ analog/dummy_l.dummy\[14\].dummy.FL analog/dummy_l.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.FL
+ analog/dummy_l.dummy\[14\].dummy.FL analog/dummy_l.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.FL
+ analog/dummy_l.dummy\[14\].dummy.FL analog/dummy_l.dummy\[14\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[14\].dummy.VREF
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[14\].dummy.VSH
+ analog/dummy_l.dummy\[14\].dummy.VREF analog/dummy_l.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[14\].dummy.VSH
+ analog/dummy_l.dummy\[14\].dummy.VREF analog/dummy_l.dummy\[14\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[14\].dummy.VREF
+ analog/dummy_l.dummy\[14\].dummy.VSH analog/dummy_l.dummy\[14\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[15\].dummy.VSH
+ analog/dummy_l.dummy\[15\].dummy.VOUTH analog/dummy_l.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[15\].dummy.VOUTH
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[15\].dummy.VOUTH
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[15\].dummy.VSH
+ analog/dummy_l.dummy\[15\].dummy.VOUTH analog/dummy_l.dummy\[15\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[15\].dummy.VSH
+ analog/dummy_l.dummy\[15\].dummy.VOUTL analog/dummy_l.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[15\].dummy.VOUTL
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[15\].dummy.VOUTL
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[15\].dummy.VSH
+ analog/dummy_l.dummy\[15\].dummy.VOUTL analog/dummy_l.dummy\[15\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.FL
+ analog/dummy_l.dummy\[15\].dummy.FL analog/dummy_l.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.FL
+ analog/dummy_l.dummy\[15\].dummy.FL analog/dummy_l.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.FL
+ analog/dummy_l.dummy\[15\].dummy.FL analog/dummy_l.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.FL
+ analog/dummy_l.dummy\[15\].dummy.FL analog/dummy_l.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.FL
+ analog/dummy_l.dummy\[15\].dummy.FL analog/dummy_l.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.FL
+ analog/dummy_l.dummy\[15\].dummy.FL analog/dummy_l.dummy\[15\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[15\].dummy.VREF
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[15\].dummy.VSH
+ analog/dummy_l.dummy\[15\].dummy.VREF analog/dummy_l.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[15\].dummy.VSH
+ analog/dummy_l.dummy\[15\].dummy.VREF analog/dummy_l.dummy\[15\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[15\].dummy.VREF
+ analog/dummy_l.dummy\[15\].dummy.VSH analog/dummy_l.dummy\[15\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[16\].dummy.VSH
+ analog/dummy_l.dummy\[16\].dummy.VOUTH analog/dummy_l.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[16\].dummy.VOUTH
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[16\].dummy.VOUTH
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[16\].dummy.VSH
+ analog/dummy_l.dummy\[16\].dummy.VOUTH analog/dummy_l.dummy\[16\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[16\].dummy.VSH
+ analog/dummy_l.dummy\[16\].dummy.VOUTL analog/dummy_l.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[16\].dummy.VOUTL
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[16\].dummy.VOUTL
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[16\].dummy.VSH
+ analog/dummy_l.dummy\[16\].dummy.VOUTL analog/dummy_l.dummy\[16\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.FL
+ analog/dummy_l.dummy\[16\].dummy.FL analog/dummy_l.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.FL
+ analog/dummy_l.dummy\[16\].dummy.FL analog/dummy_l.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.FL
+ analog/dummy_l.dummy\[16\].dummy.FL analog/dummy_l.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.FL
+ analog/dummy_l.dummy\[16\].dummy.FL analog/dummy_l.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.FL
+ analog/dummy_l.dummy\[16\].dummy.FL analog/dummy_l.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.FL
+ analog/dummy_l.dummy\[16\].dummy.FL analog/dummy_l.dummy\[16\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[16\].dummy.VREF
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[16\].dummy.VSH
+ analog/dummy_l.dummy\[16\].dummy.VREF analog/dummy_l.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[16\].dummy.VSH
+ analog/dummy_l.dummy\[16\].dummy.VREF analog/dummy_l.dummy\[16\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[16\].dummy.VREF
+ analog/dummy_l.dummy\[16\].dummy.VSH analog/dummy_l.dummy\[16\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[17\].dummy.VSH
+ analog/dummy_l.dummy\[17\].dummy.VOUTH analog/dummy_l.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[17\].dummy.VOUTH
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[17\].dummy.VOUTH
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[17\].dummy.VSH
+ analog/dummy_l.dummy\[17\].dummy.VOUTH analog/dummy_l.dummy\[17\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[17\].dummy.VSH
+ analog/dummy_l.dummy\[17\].dummy.VOUTL analog/dummy_l.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[17\].dummy.VOUTL
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[17\].dummy.VOUTL
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[17\].dummy.VSH
+ analog/dummy_l.dummy\[17\].dummy.VOUTL analog/dummy_l.dummy\[17\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.FL
+ analog/dummy_l.dummy\[17\].dummy.FL analog/dummy_l.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.FL
+ analog/dummy_l.dummy\[17\].dummy.FL analog/dummy_l.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.FL
+ analog/dummy_l.dummy\[17\].dummy.FL analog/dummy_l.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.FL
+ analog/dummy_l.dummy\[17\].dummy.FL analog/dummy_l.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.FL
+ analog/dummy_l.dummy\[17\].dummy.FL analog/dummy_l.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.FL
+ analog/dummy_l.dummy\[17\].dummy.FL analog/dummy_l.dummy\[17\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[17\].dummy.VREF
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[17\].dummy.VSH
+ analog/dummy_l.dummy\[17\].dummy.VREF analog/dummy_l.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[17\].dummy.VSH
+ analog/dummy_l.dummy\[17\].dummy.VREF analog/dummy_l.dummy\[17\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[17\].dummy.VREF
+ analog/dummy_l.dummy\[17\].dummy.VSH analog/dummy_l.dummy\[17\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[18\].dummy.VSH
+ analog/dummy_l.dummy\[18\].dummy.VOUTH analog/dummy_l.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[18\].dummy.VOUTH
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[18\].dummy.VOUTH
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[18\].dummy.VSH
+ analog/dummy_l.dummy\[18\].dummy.VOUTH analog/dummy_l.dummy\[18\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[18\].dummy.VSH
+ analog/dummy_l.dummy\[18\].dummy.VOUTL analog/dummy_l.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[18\].dummy.VOUTL
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[18\].dummy.VOUTL
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[18\].dummy.VSH
+ analog/dummy_l.dummy\[18\].dummy.VOUTL analog/dummy_l.dummy\[18\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.FL
+ analog/dummy_l.dummy\[18\].dummy.FL analog/dummy_l.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.FL
+ analog/dummy_l.dummy\[18\].dummy.FL analog/dummy_l.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.FL
+ analog/dummy_l.dummy\[18\].dummy.FL analog/dummy_l.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.FL
+ analog/dummy_l.dummy\[18\].dummy.FL analog/dummy_l.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.FL
+ analog/dummy_l.dummy\[18\].dummy.FL analog/dummy_l.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.FL
+ analog/dummy_l.dummy\[18\].dummy.FL analog/dummy_l.dummy\[18\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[18\].dummy.VREF
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[18\].dummy.VSH
+ analog/dummy_l.dummy\[18\].dummy.VREF analog/dummy_l.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[18\].dummy.VSH
+ analog/dummy_l.dummy\[18\].dummy.VREF analog/dummy_l.dummy\[18\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[18\].dummy.VREF
+ analog/dummy_l.dummy\[18\].dummy.VSH analog/dummy_l.dummy\[18\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[19\].dummy.VSH
+ analog/dummy_l.dummy\[19\].dummy.VOUTH analog/dummy_l.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[19\].dummy.VOUTH
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[19\].dummy.VOUTH
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[19\].dummy.VSH
+ analog/dummy_l.dummy\[19\].dummy.VOUTH analog/dummy_l.dummy\[19\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[19\].dummy.VSH
+ analog/dummy_l.dummy\[19\].dummy.VOUTL analog/dummy_l.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[19\].dummy.VOUTL
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[19\].dummy.VOUTL
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[19\].dummy.VSH
+ analog/dummy_l.dummy\[19\].dummy.VOUTL analog/dummy_l.dummy\[19\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.FL
+ analog/dummy_l.dummy\[19\].dummy.FL analog/dummy_l.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.FL
+ analog/dummy_l.dummy\[19\].dummy.FL analog/dummy_l.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.FL
+ analog/dummy_l.dummy\[19\].dummy.FL analog/dummy_l.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.FL
+ analog/dummy_l.dummy\[19\].dummy.FL analog/dummy_l.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.FL
+ analog/dummy_l.dummy\[19\].dummy.FL analog/dummy_l.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.FL
+ analog/dummy_l.dummy\[19\].dummy.FL analog/dummy_l.dummy\[19\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[19\].dummy.VREF
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[19\].dummy.VSH
+ analog/dummy_l.dummy\[19\].dummy.VREF analog/dummy_l.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[19\].dummy.VSH
+ analog/dummy_l.dummy\[19\].dummy.VREF analog/dummy_l.dummy\[19\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[19\].dummy.VREF
+ analog/dummy_l.dummy\[19\].dummy.VSH analog/dummy_l.dummy\[19\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[1\].dummy.VSH
+ analog/dummy_l.dummy\[1\].dummy.VOUTH analog/dummy_l.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[1\].dummy.VOUTH
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[1\].dummy.VOUTH
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[1\].dummy.VSH
+ analog/dummy_l.dummy\[1\].dummy.VOUTH analog/dummy_l.dummy\[1\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[1\].dummy.VSH
+ analog/dummy_l.dummy\[1\].dummy.VOUTL analog/dummy_l.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[1\].dummy.VOUTL
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[1\].dummy.VOUTL
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[1\].dummy.VSH
+ analog/dummy_l.dummy\[1\].dummy.VOUTL analog/dummy_l.dummy\[1\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.FL
+ analog/dummy_l.dummy\[1\].dummy.FL analog/dummy_l.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.FL
+ analog/dummy_l.dummy\[1\].dummy.FL analog/dummy_l.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.FL
+ analog/dummy_l.dummy\[1\].dummy.FL analog/dummy_l.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.FL
+ analog/dummy_l.dummy\[1\].dummy.FL analog/dummy_l.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.FL
+ analog/dummy_l.dummy\[1\].dummy.FL analog/dummy_l.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.FL
+ analog/dummy_l.dummy\[1\].dummy.FL analog/dummy_l.dummy\[1\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[1\].dummy.VREF
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[1\].dummy.VSH
+ analog/dummy_l.dummy\[1\].dummy.VREF analog/dummy_l.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[1\].dummy.VSH
+ analog/dummy_l.dummy\[1\].dummy.VREF analog/dummy_l.dummy\[1\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[1\].dummy.VREF
+ analog/dummy_l.dummy\[1\].dummy.VSH analog/dummy_l.dummy\[1\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[20\].dummy.VSH
+ analog/dummy_l.dummy\[20\].dummy.VOUTH analog/dummy_l.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[20\].dummy.VOUTH
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[20\].dummy.VOUTH
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[20\].dummy.VSH
+ analog/dummy_l.dummy\[20\].dummy.VOUTH analog/dummy_l.dummy\[20\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[20\].dummy.VSH
+ analog/dummy_l.dummy\[20\].dummy.VOUTL analog/dummy_l.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[20\].dummy.VOUTL
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[20\].dummy.VOUTL
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[20\].dummy.VSH
+ analog/dummy_l.dummy\[20\].dummy.VOUTL analog/dummy_l.dummy\[20\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.FL
+ analog/dummy_l.dummy\[20\].dummy.FL analog/dummy_l.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.FL
+ analog/dummy_l.dummy\[20\].dummy.FL analog/dummy_l.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.FL
+ analog/dummy_l.dummy\[20\].dummy.FL analog/dummy_l.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.FL
+ analog/dummy_l.dummy\[20\].dummy.FL analog/dummy_l.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.FL
+ analog/dummy_l.dummy\[20\].dummy.FL analog/dummy_l.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.FL
+ analog/dummy_l.dummy\[20\].dummy.FL analog/dummy_l.dummy\[20\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[20\].dummy.VREF
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[20\].dummy.VSH
+ analog/dummy_l.dummy\[20\].dummy.VREF analog/dummy_l.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[20\].dummy.VSH
+ analog/dummy_l.dummy\[20\].dummy.VREF analog/dummy_l.dummy\[20\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[20\].dummy.VREF
+ analog/dummy_l.dummy\[20\].dummy.VSH analog/dummy_l.dummy\[20\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[21\].dummy.VSH
+ analog/dummy_l.dummy\[21\].dummy.VOUTH analog/dummy_l.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[21\].dummy.VOUTH
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[21\].dummy.VOUTH
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[21\].dummy.VSH
+ analog/dummy_l.dummy\[21\].dummy.VOUTH analog/dummy_l.dummy\[21\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[21\].dummy.VSH
+ analog/dummy_l.dummy\[21\].dummy.VOUTL analog/dummy_l.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[21\].dummy.VOUTL
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[21\].dummy.VOUTL
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[21\].dummy.VSH
+ analog/dummy_l.dummy\[21\].dummy.VOUTL analog/dummy_l.dummy\[21\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.FL
+ analog/dummy_l.dummy\[21\].dummy.FL analog/dummy_l.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.FL
+ analog/dummy_l.dummy\[21\].dummy.FL analog/dummy_l.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.FL
+ analog/dummy_l.dummy\[21\].dummy.FL analog/dummy_l.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.FL
+ analog/dummy_l.dummy\[21\].dummy.FL analog/dummy_l.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.FL
+ analog/dummy_l.dummy\[21\].dummy.FL analog/dummy_l.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.FL
+ analog/dummy_l.dummy\[21\].dummy.FL analog/dummy_l.dummy\[21\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[21\].dummy.VREF
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[21\].dummy.VSH
+ analog/dummy_l.dummy\[21\].dummy.VREF analog/dummy_l.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[21\].dummy.VSH
+ analog/dummy_l.dummy\[21\].dummy.VREF analog/dummy_l.dummy\[21\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[21\].dummy.VREF
+ analog/dummy_l.dummy\[21\].dummy.VSH analog/dummy_l.dummy\[21\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[22\].dummy.VSH
+ analog/dummy_l.dummy\[22\].dummy.VOUTH analog/dummy_l.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[22\].dummy.VOUTH
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[22\].dummy.VOUTH
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[22\].dummy.VSH
+ analog/dummy_l.dummy\[22\].dummy.VOUTH analog/dummy_l.dummy\[22\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[22\].dummy.VSH
+ analog/dummy_l.dummy\[22\].dummy.VOUTL analog/dummy_l.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[22\].dummy.VOUTL
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[22\].dummy.VOUTL
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[22\].dummy.VSH
+ analog/dummy_l.dummy\[22\].dummy.VOUTL analog/dummy_l.dummy\[22\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.FL
+ analog/dummy_l.dummy\[22\].dummy.FL analog/dummy_l.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.FL
+ analog/dummy_l.dummy\[22\].dummy.FL analog/dummy_l.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.FL
+ analog/dummy_l.dummy\[22\].dummy.FL analog/dummy_l.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.FL
+ analog/dummy_l.dummy\[22\].dummy.FL analog/dummy_l.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.FL
+ analog/dummy_l.dummy\[22\].dummy.FL analog/dummy_l.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.FL
+ analog/dummy_l.dummy\[22\].dummy.FL analog/dummy_l.dummy\[22\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[22\].dummy.VREF
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[22\].dummy.VSH
+ analog/dummy_l.dummy\[22\].dummy.VREF analog/dummy_l.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[22\].dummy.VSH
+ analog/dummy_l.dummy\[22\].dummy.VREF analog/dummy_l.dummy\[22\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[22\].dummy.VREF
+ analog/dummy_l.dummy\[22\].dummy.VSH analog/dummy_l.dummy\[22\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[23\].dummy.VSH
+ analog/dummy_l.dummy\[23\].dummy.VOUTH analog/dummy_l.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[23\].dummy.VOUTH
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[23\].dummy.VOUTH
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[23\].dummy.VSH
+ analog/dummy_l.dummy\[23\].dummy.VOUTH analog/dummy_l.dummy\[23\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[23\].dummy.VSH
+ analog/dummy_l.dummy\[23\].dummy.VOUTL analog/dummy_l.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[23\].dummy.VOUTL
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[23\].dummy.VOUTL
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[23\].dummy.VSH
+ analog/dummy_l.dummy\[23\].dummy.VOUTL analog/dummy_l.dummy\[23\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.FL
+ analog/dummy_l.dummy\[23\].dummy.FL analog/dummy_l.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.FL
+ analog/dummy_l.dummy\[23\].dummy.FL analog/dummy_l.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.FL
+ analog/dummy_l.dummy\[23\].dummy.FL analog/dummy_l.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.FL
+ analog/dummy_l.dummy\[23\].dummy.FL analog/dummy_l.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.FL
+ analog/dummy_l.dummy\[23\].dummy.FL analog/dummy_l.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.FL
+ analog/dummy_l.dummy\[23\].dummy.FL analog/dummy_l.dummy\[23\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[23\].dummy.VREF
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[23\].dummy.VSH
+ analog/dummy_l.dummy\[23\].dummy.VREF analog/dummy_l.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[23\].dummy.VSH
+ analog/dummy_l.dummy\[23\].dummy.VREF analog/dummy_l.dummy\[23\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[23\].dummy.VREF
+ analog/dummy_l.dummy\[23\].dummy.VSH analog/dummy_l.dummy\[23\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[24\].dummy.VSH
+ analog/dummy_l.dummy\[24\].dummy.VOUTH analog/dummy_l.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[24\].dummy.VOUTH
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[24\].dummy.VOUTH
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[24\].dummy.VSH
+ analog/dummy_l.dummy\[24\].dummy.VOUTH analog/dummy_l.dummy\[24\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[24\].dummy.VSH
+ analog/dummy_l.dummy\[24\].dummy.VOUTL analog/dummy_l.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[24\].dummy.VOUTL
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[24\].dummy.VOUTL
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[24\].dummy.VSH
+ analog/dummy_l.dummy\[24\].dummy.VOUTL analog/dummy_l.dummy\[24\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.FL
+ analog/dummy_l.dummy\[24\].dummy.FL analog/dummy_l.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.FL
+ analog/dummy_l.dummy\[24\].dummy.FL analog/dummy_l.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.FL
+ analog/dummy_l.dummy\[24\].dummy.FL analog/dummy_l.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.FL
+ analog/dummy_l.dummy\[24\].dummy.FL analog/dummy_l.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.FL
+ analog/dummy_l.dummy\[24\].dummy.FL analog/dummy_l.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.FL
+ analog/dummy_l.dummy\[24\].dummy.FL analog/dummy_l.dummy\[24\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[24\].dummy.VREF
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[24\].dummy.VSH
+ analog/dummy_l.dummy\[24\].dummy.VREF analog/dummy_l.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[24\].dummy.VSH
+ analog/dummy_l.dummy\[24\].dummy.VREF analog/dummy_l.dummy\[24\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[24\].dummy.VREF
+ analog/dummy_l.dummy\[24\].dummy.VSH analog/dummy_l.dummy\[24\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[25\].dummy.VSH
+ analog/dummy_l.dummy\[25\].dummy.VOUTH analog/dummy_l.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[25\].dummy.VOUTH
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[25\].dummy.VOUTH
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[25\].dummy.VSH
+ analog/dummy_l.dummy\[25\].dummy.VOUTH analog/dummy_l.dummy\[25\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[25\].dummy.VSH
+ analog/dummy_l.dummy\[25\].dummy.VOUTL analog/dummy_l.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[25\].dummy.VOUTL
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[25\].dummy.VOUTL
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[25\].dummy.VSH
+ analog/dummy_l.dummy\[25\].dummy.VOUTL analog/dummy_l.dummy\[25\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.FL
+ analog/dummy_l.dummy\[25\].dummy.FL analog/dummy_l.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.FL
+ analog/dummy_l.dummy\[25\].dummy.FL analog/dummy_l.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.FL
+ analog/dummy_l.dummy\[25\].dummy.FL analog/dummy_l.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.FL
+ analog/dummy_l.dummy\[25\].dummy.FL analog/dummy_l.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.FL
+ analog/dummy_l.dummy\[25\].dummy.FL analog/dummy_l.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.FL
+ analog/dummy_l.dummy\[25\].dummy.FL analog/dummy_l.dummy\[25\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[25\].dummy.VREF
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[25\].dummy.VSH
+ analog/dummy_l.dummy\[25\].dummy.VREF analog/dummy_l.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[25\].dummy.VSH
+ analog/dummy_l.dummy\[25\].dummy.VREF analog/dummy_l.dummy\[25\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[25\].dummy.VREF
+ analog/dummy_l.dummy\[25\].dummy.VSH analog/dummy_l.dummy\[25\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[26\].dummy.VSH
+ analog/dummy_l.dummy\[26\].dummy.VOUTH analog/dummy_l.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[26\].dummy.VOUTH
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[26\].dummy.VOUTH
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[26\].dummy.VSH
+ analog/dummy_l.dummy\[26\].dummy.VOUTH analog/dummy_l.dummy\[26\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[26\].dummy.VSH
+ analog/dummy_l.dummy\[26\].dummy.VOUTL analog/dummy_l.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[26\].dummy.VOUTL
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[26\].dummy.VOUTL
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[26\].dummy.VSH
+ analog/dummy_l.dummy\[26\].dummy.VOUTL analog/dummy_l.dummy\[26\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.FL
+ analog/dummy_l.dummy\[26\].dummy.FL analog/dummy_l.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.FL
+ analog/dummy_l.dummy\[26\].dummy.FL analog/dummy_l.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.FL
+ analog/dummy_l.dummy\[26\].dummy.FL analog/dummy_l.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.FL
+ analog/dummy_l.dummy\[26\].dummy.FL analog/dummy_l.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.FL
+ analog/dummy_l.dummy\[26\].dummy.FL analog/dummy_l.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.FL
+ analog/dummy_l.dummy\[26\].dummy.FL analog/dummy_l.dummy\[26\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[26\].dummy.VREF
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[26\].dummy.VSH
+ analog/dummy_l.dummy\[26\].dummy.VREF analog/dummy_l.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[26\].dummy.VSH
+ analog/dummy_l.dummy\[26\].dummy.VREF analog/dummy_l.dummy\[26\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[26\].dummy.VREF
+ analog/dummy_l.dummy\[26\].dummy.VSH analog/dummy_l.dummy\[26\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[27\].dummy.VSH
+ analog/dummy_l.dummy\[27\].dummy.VOUTH analog/dummy_l.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[27\].dummy.VOUTH
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[27\].dummy.VOUTH
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[27\].dummy.VSH
+ analog/dummy_l.dummy\[27\].dummy.VOUTH analog/dummy_l.dummy\[27\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[27\].dummy.VSH
+ analog/dummy_l.dummy\[27\].dummy.VOUTL analog/dummy_l.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[27\].dummy.VOUTL
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[27\].dummy.VOUTL
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[27\].dummy.VSH
+ analog/dummy_l.dummy\[27\].dummy.VOUTL analog/dummy_l.dummy\[27\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.FL
+ analog/dummy_l.dummy\[27\].dummy.FL analog/dummy_l.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.FL
+ analog/dummy_l.dummy\[27\].dummy.FL analog/dummy_l.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.FL
+ analog/dummy_l.dummy\[27\].dummy.FL analog/dummy_l.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.FL
+ analog/dummy_l.dummy\[27\].dummy.FL analog/dummy_l.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.FL
+ analog/dummy_l.dummy\[27\].dummy.FL analog/dummy_l.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.FL
+ analog/dummy_l.dummy\[27\].dummy.FL analog/dummy_l.dummy\[27\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[27\].dummy.VREF
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[27\].dummy.VSH
+ analog/dummy_l.dummy\[27\].dummy.VREF analog/dummy_l.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[27\].dummy.VSH
+ analog/dummy_l.dummy\[27\].dummy.VREF analog/dummy_l.dummy\[27\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[27\].dummy.VREF
+ analog/dummy_l.dummy\[27\].dummy.VSH analog/dummy_l.dummy\[27\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[2\].dummy.VSH
+ analog/dummy_l.dummy\[2\].dummy.VOUTH analog/dummy_l.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[2\].dummy.VOUTH
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[2\].dummy.VOUTH
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[2\].dummy.VSH
+ analog/dummy_l.dummy\[2\].dummy.VOUTH analog/dummy_l.dummy\[2\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[2\].dummy.VSH
+ analog/dummy_l.dummy\[2\].dummy.VOUTL analog/dummy_l.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[2\].dummy.VOUTL
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[2\].dummy.VOUTL
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[2\].dummy.VSH
+ analog/dummy_l.dummy\[2\].dummy.VOUTL analog/dummy_l.dummy\[2\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.FL
+ analog/dummy_l.dummy\[2\].dummy.FL analog/dummy_l.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.FL
+ analog/dummy_l.dummy\[2\].dummy.FL analog/dummy_l.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.FL
+ analog/dummy_l.dummy\[2\].dummy.FL analog/dummy_l.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.FL
+ analog/dummy_l.dummy\[2\].dummy.FL analog/dummy_l.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.FL
+ analog/dummy_l.dummy\[2\].dummy.FL analog/dummy_l.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.FL
+ analog/dummy_l.dummy\[2\].dummy.FL analog/dummy_l.dummy\[2\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[2\].dummy.VREF
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[2\].dummy.VSH
+ analog/dummy_l.dummy\[2\].dummy.VREF analog/dummy_l.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[2\].dummy.VSH
+ analog/dummy_l.dummy\[2\].dummy.VREF analog/dummy_l.dummy\[2\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[2\].dummy.VREF
+ analog/dummy_l.dummy\[2\].dummy.VSH analog/dummy_l.dummy\[2\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[3\].dummy.VSH
+ analog/dummy_l.dummy\[3\].dummy.VOUTH analog/dummy_l.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[3\].dummy.VOUTH
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[3\].dummy.VOUTH
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[3\].dummy.VSH
+ analog/dummy_l.dummy\[3\].dummy.VOUTH analog/dummy_l.dummy\[3\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[3\].dummy.VSH
+ analog/dummy_l.dummy\[3\].dummy.VOUTL analog/dummy_l.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[3\].dummy.VOUTL
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[3\].dummy.VOUTL
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[3\].dummy.VSH
+ analog/dummy_l.dummy\[3\].dummy.VOUTL analog/dummy_l.dummy\[3\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.FL
+ analog/dummy_l.dummy\[3\].dummy.FL analog/dummy_l.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.FL
+ analog/dummy_l.dummy\[3\].dummy.FL analog/dummy_l.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.FL
+ analog/dummy_l.dummy\[3\].dummy.FL analog/dummy_l.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.FL
+ analog/dummy_l.dummy\[3\].dummy.FL analog/dummy_l.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.FL
+ analog/dummy_l.dummy\[3\].dummy.FL analog/dummy_l.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.FL
+ analog/dummy_l.dummy\[3\].dummy.FL analog/dummy_l.dummy\[3\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[3\].dummy.VREF
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[3\].dummy.VSH
+ analog/dummy_l.dummy\[3\].dummy.VREF analog/dummy_l.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[3\].dummy.VSH
+ analog/dummy_l.dummy\[3\].dummy.VREF analog/dummy_l.dummy\[3\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[3\].dummy.VREF
+ analog/dummy_l.dummy\[3\].dummy.VSH analog/dummy_l.dummy\[3\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[4\].dummy.VSH
+ analog/dummy_l.dummy\[4\].dummy.VOUTH analog/dummy_l.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[4\].dummy.VOUTH
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[4\].dummy.VOUTH
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[4\].dummy.VSH
+ analog/dummy_l.dummy\[4\].dummy.VOUTH analog/dummy_l.dummy\[4\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[4\].dummy.VSH
+ analog/dummy_l.dummy\[4\].dummy.VOUTL analog/dummy_l.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[4\].dummy.VOUTL
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[4\].dummy.VOUTL
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[4\].dummy.VSH
+ analog/dummy_l.dummy\[4\].dummy.VOUTL analog/dummy_l.dummy\[4\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.FL
+ analog/dummy_l.dummy\[4\].dummy.FL analog/dummy_l.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.FL
+ analog/dummy_l.dummy\[4\].dummy.FL analog/dummy_l.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.FL
+ analog/dummy_l.dummy\[4\].dummy.FL analog/dummy_l.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.FL
+ analog/dummy_l.dummy\[4\].dummy.FL analog/dummy_l.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.FL
+ analog/dummy_l.dummy\[4\].dummy.FL analog/dummy_l.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.FL
+ analog/dummy_l.dummy\[4\].dummy.FL analog/dummy_l.dummy\[4\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[4\].dummy.VREF
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[4\].dummy.VSH
+ analog/dummy_l.dummy\[4\].dummy.VREF analog/dummy_l.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[4\].dummy.VSH
+ analog/dummy_l.dummy\[4\].dummy.VREF analog/dummy_l.dummy\[4\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[4\].dummy.VREF
+ analog/dummy_l.dummy\[4\].dummy.VSH analog/dummy_l.dummy\[4\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[5\].dummy.VSH
+ analog/dummy_l.dummy\[5\].dummy.VOUTH analog/dummy_l.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[5\].dummy.VOUTH
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[5\].dummy.VOUTH
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[5\].dummy.VSH
+ analog/dummy_l.dummy\[5\].dummy.VOUTH analog/dummy_l.dummy\[5\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[5\].dummy.VSH
+ analog/dummy_l.dummy\[5\].dummy.VOUTL analog/dummy_l.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[5\].dummy.VOUTL
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[5\].dummy.VOUTL
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[5\].dummy.VSH
+ analog/dummy_l.dummy\[5\].dummy.VOUTL analog/dummy_l.dummy\[5\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.FL
+ analog/dummy_l.dummy\[5\].dummy.FL analog/dummy_l.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.FL
+ analog/dummy_l.dummy\[5\].dummy.FL analog/dummy_l.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.FL
+ analog/dummy_l.dummy\[5\].dummy.FL analog/dummy_l.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.FL
+ analog/dummy_l.dummy\[5\].dummy.FL analog/dummy_l.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.FL
+ analog/dummy_l.dummy\[5\].dummy.FL analog/dummy_l.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.FL
+ analog/dummy_l.dummy\[5\].dummy.FL analog/dummy_l.dummy\[5\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[5\].dummy.VREF
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[5\].dummy.VSH
+ analog/dummy_l.dummy\[5\].dummy.VREF analog/dummy_l.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[5\].dummy.VSH
+ analog/dummy_l.dummy\[5\].dummy.VREF analog/dummy_l.dummy\[5\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[5\].dummy.VREF
+ analog/dummy_l.dummy\[5\].dummy.VSH analog/dummy_l.dummy\[5\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[6\].dummy.VSH
+ analog/dummy_l.dummy\[6\].dummy.VOUTH analog/dummy_l.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[6\].dummy.VOUTH
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[6\].dummy.VOUTH
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[6\].dummy.VSH
+ analog/dummy_l.dummy\[6\].dummy.VOUTH analog/dummy_l.dummy\[6\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[6\].dummy.VSH
+ analog/dummy_l.dummy\[6\].dummy.VOUTL analog/dummy_l.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[6\].dummy.VOUTL
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[6\].dummy.VOUTL
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[6\].dummy.VSH
+ analog/dummy_l.dummy\[6\].dummy.VOUTL analog/dummy_l.dummy\[6\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.FL
+ analog/dummy_l.dummy\[6\].dummy.FL analog/dummy_l.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.FL
+ analog/dummy_l.dummy\[6\].dummy.FL analog/dummy_l.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.FL
+ analog/dummy_l.dummy\[6\].dummy.FL analog/dummy_l.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.FL
+ analog/dummy_l.dummy\[6\].dummy.FL analog/dummy_l.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.FL
+ analog/dummy_l.dummy\[6\].dummy.FL analog/dummy_l.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.FL
+ analog/dummy_l.dummy\[6\].dummy.FL analog/dummy_l.dummy\[6\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[6\].dummy.VREF
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[6\].dummy.VSH
+ analog/dummy_l.dummy\[6\].dummy.VREF analog/dummy_l.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[6\].dummy.VSH
+ analog/dummy_l.dummy\[6\].dummy.VREF analog/dummy_l.dummy\[6\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[6\].dummy.VREF
+ analog/dummy_l.dummy\[6\].dummy.VSH analog/dummy_l.dummy\[6\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[7\].dummy.VSH
+ analog/dummy_l.dummy\[7\].dummy.VOUTH analog/dummy_l.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[7\].dummy.VOUTH
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[7\].dummy.VOUTH
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[7\].dummy.VSH
+ analog/dummy_l.dummy\[7\].dummy.VOUTH analog/dummy_l.dummy\[7\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[7\].dummy.VSH
+ analog/dummy_l.dummy\[7\].dummy.VOUTL analog/dummy_l.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[7\].dummy.VOUTL
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[7\].dummy.VOUTL
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[7\].dummy.VSH
+ analog/dummy_l.dummy\[7\].dummy.VOUTL analog/dummy_l.dummy\[7\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.FL
+ analog/dummy_l.dummy\[7\].dummy.FL analog/dummy_l.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.FL
+ analog/dummy_l.dummy\[7\].dummy.FL analog/dummy_l.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.FL
+ analog/dummy_l.dummy\[7\].dummy.FL analog/dummy_l.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.FL
+ analog/dummy_l.dummy\[7\].dummy.FL analog/dummy_l.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.FL
+ analog/dummy_l.dummy\[7\].dummy.FL analog/dummy_l.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.FL
+ analog/dummy_l.dummy\[7\].dummy.FL analog/dummy_l.dummy\[7\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[7\].dummy.VREF
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[7\].dummy.VSH
+ analog/dummy_l.dummy\[7\].dummy.VREF analog/dummy_l.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[7\].dummy.VSH
+ analog/dummy_l.dummy\[7\].dummy.VREF analog/dummy_l.dummy\[7\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[7\].dummy.VREF
+ analog/dummy_l.dummy\[7\].dummy.VSH analog/dummy_l.dummy\[7\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[8\].dummy.VSH
+ analog/dummy_l.dummy\[8\].dummy.VOUTH analog/dummy_l.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[8\].dummy.VOUTH
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[8\].dummy.VOUTH
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[8\].dummy.VSH
+ analog/dummy_l.dummy\[8\].dummy.VOUTH analog/dummy_l.dummy\[8\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[8\].dummy.VSH
+ analog/dummy_l.dummy\[8\].dummy.VOUTL analog/dummy_l.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[8\].dummy.VOUTL
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[8\].dummy.VOUTL
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[8\].dummy.VSH
+ analog/dummy_l.dummy\[8\].dummy.VOUTL analog/dummy_l.dummy\[8\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.FL
+ analog/dummy_l.dummy\[8\].dummy.FL analog/dummy_l.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.FL
+ analog/dummy_l.dummy\[8\].dummy.FL analog/dummy_l.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.FL
+ analog/dummy_l.dummy\[8\].dummy.FL analog/dummy_l.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.FL
+ analog/dummy_l.dummy\[8\].dummy.FL analog/dummy_l.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.FL
+ analog/dummy_l.dummy\[8\].dummy.FL analog/dummy_l.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.FL
+ analog/dummy_l.dummy\[8\].dummy.FL analog/dummy_l.dummy\[8\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[8\].dummy.VREF
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[8\].dummy.VSH
+ analog/dummy_l.dummy\[8\].dummy.VREF analog/dummy_l.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[8\].dummy.VSH
+ analog/dummy_l.dummy\[8\].dummy.VREF analog/dummy_l.dummy\[8\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[8\].dummy.VREF
+ analog/dummy_l.dummy\[8\].dummy.VSH analog/dummy_l.dummy\[8\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[9\].dummy.VSH
+ analog/dummy_l.dummy\[9\].dummy.VOUTH analog/dummy_l.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[9\].dummy.VOUTH
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[9\].dummy.VOUTH
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[9\].dummy.VSH
+ analog/dummy_l.dummy\[9\].dummy.VOUTH analog/dummy_l.dummy\[9\].dummy.VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[9\].dummy.VSH
+ analog/dummy_l.dummy\[9\].dummy.VOUTL analog/dummy_l.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[9\].dummy.VOUTL
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[9\].dummy.VOUTL
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[9\].dummy.VSH
+ analog/dummy_l.dummy\[9\].dummy.VOUTL analog/dummy_l.dummy\[9\].dummy.VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap\[0\].cap/impl
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.FL
+ analog/dummy_l.dummy\[9\].dummy.FL analog/dummy_l.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap\[1\].cap/impl
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.FL
+ analog/dummy_l.dummy\[9\].dummy.FL analog/dummy_l.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap\[2\].cap/impl
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.FL
+ analog/dummy_l.dummy\[9\].dummy.FL analog/dummy_l.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap\[3\].cap/impl
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.FL
+ analog/dummy_l.dummy\[9\].dummy.FL analog/dummy_l.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap\[4\].cap/impl
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.FL
+ analog/dummy_l.dummy\[9\].dummy.FL analog/dummy_l.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap\[5\].cap/impl
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.FL
+ analog/dummy_l.dummy\[9\].dummy.FL analog/dummy_l.dummy\[9\].dummy.FL
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[9\].dummy.VREF
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRH analog/dummy_l.dummy\[9\].dummy.VSH
+ analog/dummy_l.dummy\[9\].dummy.VREF analog/dummy_l.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[9\].dummy.VSH
+ analog/dummy_l.dummy\[9\].dummy.VREF analog/dummy_l.dummy\[9\].dummy.VREF
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/dummy_l.dummy\[0\].dummy.CRHB analog/dummy_l.dummy\[9\].dummy.VREF
+ analog/dummy_l.dummy\[9\].dummy.VSH analog/dummy_l.dummy\[9\].dummy.VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/dummy_l.tieh.impl AVDD VSS analog/dummy_l.dummy\[0\].dummy.CRHB
+ sg13g2f_TIEH
Xanalog/dummy_l.tiel.impl AVDD VSS analog/dummy_l.dummy\[0\].dummy.CRH
+ sg13g2f_TIEL
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[0\] analog/LSB_H_VSH\[1\] analog/VOUTH analog/LSB_H_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[0\] analog/VOUTH analog/LSB_H_VSH\[1\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[0\] analog/VOUTH analog/LSB_H_VSH\[1\] analog/LSB_H_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[0\] analog/LSB_H_VSH\[1\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[0\] analog/LSB_H_VSH\[1\] analog/VOUTL analog/LSB_H_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[0\] analog/VOUTL analog/LSB_H_VSH\[1\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[0\] analog/VOUTL analog/LSB_H_VSH\[1\] analog/LSB_H_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[0\] analog/LSB_H_VSH\[1\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap\[0\].cap/impl
+ analog/LSB_H_VSH\[1\] analog/LSB_H_FL\[1\] analog/LSB_H_FL\[1\]
+ analog/LSB_H_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap\[1\].cap/impl
+ analog/LSB_H_VSH\[1\] analog/LSB_H_FL\[1\] analog/LSB_H_FL\[1\]
+ analog/LSB_H_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap\[2\].cap/impl
+ analog/LSB_H_VSH\[1\] analog/LSB_H_FL\[1\] analog/LSB_H_FL\[1\]
+ analog/LSB_H_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap\[3\].cap/impl
+ analog/LSB_H_VSH\[1\] analog/LSB_H_FL\[1\] analog/LSB_H_FL\[1\]
+ analog/LSB_H_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap\[4\].cap/impl
+ analog/LSB_H_VSH\[1\] analog/LSB_H_FL\[1\] analog/LSB_H_FL\[1\]
+ analog/LSB_H_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap\[5\].cap/impl
+ analog/LSB_H_VSH\[1\] analog/LSB_H_FL\[1\] analog/LSB_H_FL\[1\]
+ analog/LSB_H_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[1\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[1\] VREFH analog/LSB_H_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[1\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[1\] analog/LSB_H_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[1\] analog/LSB_H_VSH\[2\] analog/VOUTH analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[1\] analog/VOUTH analog/LSB_H_VSH\[2\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[1\] analog/VOUTH analog/LSB_H_VSH\[2\] analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[1\] analog/LSB_H_VSH\[2\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[1\] analog/LSB_H_VSH\[2\] analog/VOUTH analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[1\] analog/VOUTH analog/LSB_H_VSH\[2\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[1\] analog/VOUTH analog/LSB_H_VSH\[2\] analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[1\] analog/LSB_H_VSH\[2\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[1\] analog/LSB_H_VSH\[2\] analog/VOUTL analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[1\] analog/VOUTL analog/LSB_H_VSH\[2\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[1\] analog/VOUTL analog/LSB_H_VSH\[2\] analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[1\] analog/LSB_H_VSH\[2\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[1\] analog/LSB_H_VSH\[2\] analog/VOUTL analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[1\] analog/VOUTL analog/LSB_H_VSH\[2\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[1\] analog/VOUTL analog/LSB_H_VSH\[2\] analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[1\] analog/LSB_H_VSH\[2\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[0\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[10\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[11\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[1\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[2\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[3\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[4\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[5\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[6\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[7\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[8\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap\[9\].cap/impl
+ analog/LSB_H_VSH\[2\] analog/LSB_H_FL\[2\] analog/LSB_H_FL\[2\]
+ analog/LSB_H_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[2\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[2\] VREFH analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[2\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[2\] analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[2\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[2\] VREFH analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[2\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[2\] analog/LSB_H_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[2\] analog/LSB_H_VSH\[3\] analog/VOUTH analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[2\] analog/VOUTH analog/LSB_H_VSH\[3\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[2\] analog/VOUTH analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[2\] analog/LSB_H_VSH\[3\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[2\] analog/LSB_H_VSH\[3\] analog/VOUTH analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[2\] analog/VOUTH analog/LSB_H_VSH\[3\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[2\] analog/VOUTH analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[2\] analog/LSB_H_VSH\[3\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[2\] analog/LSB_H_VSH\[3\] analog/VOUTH analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[2\] analog/VOUTH analog/LSB_H_VSH\[3\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[2\] analog/VOUTH analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[2\] analog/LSB_H_VSH\[3\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[2\] analog/LSB_H_VSH\[3\] analog/VOUTH analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[2\] analog/VOUTH analog/LSB_H_VSH\[3\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[2\] analog/VOUTH analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[2\] analog/LSB_H_VSH\[3\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[2\] analog/LSB_H_VSH\[3\] analog/VOUTL analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[2\] analog/VOUTL analog/LSB_H_VSH\[3\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[2\] analog/VOUTL analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[2\] analog/LSB_H_VSH\[3\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[2\] analog/LSB_H_VSH\[3\] analog/VOUTL analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[2\] analog/VOUTL analog/LSB_H_VSH\[3\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[2\] analog/VOUTL analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[2\] analog/LSB_H_VSH\[3\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[2\] analog/LSB_H_VSH\[3\] analog/VOUTL analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[2\] analog/VOUTL analog/LSB_H_VSH\[3\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[2\] analog/VOUTL analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[2\] analog/LSB_H_VSH\[3\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[2\] analog/LSB_H_VSH\[3\] analog/VOUTL analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[2\] analog/VOUTL analog/LSB_H_VSH\[3\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[2\] analog/VOUTL analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[2\] analog/LSB_H_VSH\[3\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[0\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[10\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[11\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[12\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[13\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[14\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[15\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[16\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[17\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[18\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[19\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[1\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[20\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[21\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[22\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[23\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[2\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[3\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[4\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[5\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[6\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[7\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[8\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap\[9\].cap/impl
+ analog/LSB_H_VSH\[3\] analog/LSB_H_FL\[3\] analog/LSB_H_FL\[3\]
+ analog/LSB_H_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[3\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[3\] VREFH analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[3\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[3\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[3\] VREFH analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[3\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[3\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[3\] VREFH analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[3\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[3\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[3\] VREFH analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[3\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[3\] analog/LSB_H_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTL analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_H_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[0\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[10\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[11\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[12\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[13\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[14\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[15\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[16\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[17\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[18\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[19\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[1\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[20\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[21\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[22\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[23\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[24\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[25\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[26\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[27\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[28\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[29\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[2\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[30\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[31\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[32\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[33\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[34\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[35\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[36\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[37\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[38\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[39\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[3\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[40\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[41\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[42\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[43\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[44\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[45\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[46\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[47\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[4\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[5\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[6\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[7\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[8\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap\[9\].cap/impl
+ analog/LSB_H_VSH\[4\] analog/LSB_H_FL\[4\] analog/LSB_H_FL\[4\]
+ analog/LSB_H_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[4\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[4\] VREFH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[4\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[4\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[4\] VREFH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[4\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[4\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[4\] VREFH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[4\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[4\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[4\] VREFH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[4\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[4\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[4\] VREFH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[4\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[4\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[4\] VREFH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[4\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[4\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[4\] VREFH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[4\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[4\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[4\] VREFH analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[4\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[4\] analog/LSB_H_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/lsb_cdac_h.cdac_unit.CRH analog/LSB_H_VSH\[0\] analog/VOUTH
+ analog/LSB_H_VSH\[0\] AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/lsb_cdac_h.cdac_unit.CRH analog/VOUTH analog/LSB_H_VSH\[0\]
+ analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/lsb_cdac_h.cdac_unit.CRHB analog/VOUTH analog/LSB_H_VSH\[0\]
+ analog/LSB_H_VSH\[0\] AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/lsb_cdac_h.cdac_unit.CRHB analog/LSB_H_VSH\[0\] analog/VOUTH
+ analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/lsb_cdac_h.cdac_unit.CRH analog/LSB_H_VSH\[0\] analog/VOUTL
+ analog/LSB_H_VSH\[0\] AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/lsb_cdac_h.cdac_unit.CRH analog/VOUTL analog/LSB_H_VSH\[0\]
+ analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/lsb_cdac_h.cdac_unit.CRHB analog/VOUTL analog/LSB_H_VSH\[0\]
+ analog/LSB_H_VSH\[0\] AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/lsb_cdac_h.cdac_unit.CRHB analog/LSB_H_VSH\[0\] analog/VOUTL
+ analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.cap\[0\].cap/impl analog/LSB_H_VSH\[0\]
+ analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_unit.cap\[1\].cap/impl analog/LSB_H_VSH\[0\]
+ analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_unit.cap\[2\].cap/impl analog/LSB_H_VSH\[0\]
+ analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_unit.cap\[3\].cap/impl analog/LSB_H_VSH\[0\]
+ analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_unit.cap\[4\].cap/impl analog/LSB_H_VSH\[0\]
+ analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_unit.cap\[5\].cap/impl analog/LSB_H_VSH\[0\]
+ analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\] analog/LSB_H_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFH analog/LSB_H_VSH\[0\] VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_H_VSH\[0\] VREFH analog/LSB_H_VSH\[0\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_H_VSH\[0\] VREFH VREFH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFH analog/LSB_H_VSH\[0\] analog/LSB_H_VSH\[0\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_h.tieh.impl AVDD VSS analog/lsb_cdac_h.cdac_unit.CRHB
+ sg13g2f_TIEH
Xanalog/lsb_cdac_h.tiel.impl AVDD VSS analog/lsb_cdac_h.cdac_unit.CRH
+ sg13g2f_TIEL
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[0\] analog/LSB_L_VSH\[1\] analog/VOUTL analog/LSB_L_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[0\] analog/VOUTL analog/LSB_L_VSH\[1\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[0\] analog/VOUTL analog/LSB_L_VSH\[1\] analog/LSB_L_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[0\] analog/LSB_L_VSH\[1\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[0\] analog/LSB_L_VSH\[1\] analog/VOUTH analog/LSB_L_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[0\] analog/VOUTH analog/LSB_L_VSH\[1\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[0\] analog/VOUTH analog/LSB_L_VSH\[1\] analog/LSB_L_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[0\] analog/LSB_L_VSH\[1\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap\[0\].cap/impl
+ analog/LSB_L_VSH\[1\] analog/LSB_L_FL\[1\] analog/LSB_L_FL\[1\]
+ analog/LSB_L_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap\[1\].cap/impl
+ analog/LSB_L_VSH\[1\] analog/LSB_L_FL\[1\] analog/LSB_L_FL\[1\]
+ analog/LSB_L_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap\[2\].cap/impl
+ analog/LSB_L_VSH\[1\] analog/LSB_L_FL\[1\] analog/LSB_L_FL\[1\]
+ analog/LSB_L_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap\[3\].cap/impl
+ analog/LSB_L_VSH\[1\] analog/LSB_L_FL\[1\] analog/LSB_L_FL\[1\]
+ analog/LSB_L_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap\[4\].cap/impl
+ analog/LSB_L_VSH\[1\] analog/LSB_L_FL\[1\] analog/LSB_L_FL\[1\]
+ analog/LSB_L_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap\[5\].cap/impl
+ analog/LSB_L_VSH\[1\] analog/LSB_L_FL\[1\] analog/LSB_L_FL\[1\]
+ analog/LSB_L_FL\[1\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[1\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[1\] VREFL analog/LSB_L_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[1\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[1\] analog/LSB_L_VSH\[1\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[1\] analog/LSB_L_VSH\[2\] analog/VOUTL analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[1\] analog/VOUTL analog/LSB_L_VSH\[2\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[1\] analog/VOUTL analog/LSB_L_VSH\[2\] analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[1\] analog/LSB_L_VSH\[2\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[1\] analog/LSB_L_VSH\[2\] analog/VOUTL analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[1\] analog/VOUTL analog/LSB_L_VSH\[2\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[1\] analog/VOUTL analog/LSB_L_VSH\[2\] analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[1\] analog/LSB_L_VSH\[2\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[1\] analog/LSB_L_VSH\[2\] analog/VOUTH analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[1\] analog/VOUTH analog/LSB_L_VSH\[2\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[1\] analog/VOUTH analog/LSB_L_VSH\[2\] analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[1\] analog/LSB_L_VSH\[2\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[1\] analog/LSB_L_VSH\[2\] analog/VOUTH analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[1\] analog/VOUTH analog/LSB_L_VSH\[2\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[1\] analog/VOUTH analog/LSB_L_VSH\[2\] analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[1\] analog/LSB_L_VSH\[2\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[0\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[10\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[11\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[1\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[2\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[3\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[4\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[5\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[6\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[7\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[8\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap\[9\].cap/impl
+ analog/LSB_L_VSH\[2\] analog/LSB_L_FL\[2\] analog/LSB_L_FL\[2\]
+ analog/LSB_L_FL\[2\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[2\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[2\] VREFL analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[2\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[2\] analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[2\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[2\] VREFL analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[2\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[2\] analog/LSB_L_VSH\[2\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[2\] analog/LSB_L_VSH\[3\] analog/VOUTL analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[2\] analog/VOUTL analog/LSB_L_VSH\[3\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[2\] analog/VOUTL analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[2\] analog/LSB_L_VSH\[3\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[2\] analog/LSB_L_VSH\[3\] analog/VOUTL analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[2\] analog/VOUTL analog/LSB_L_VSH\[3\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[2\] analog/VOUTL analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[2\] analog/LSB_L_VSH\[3\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[2\] analog/LSB_L_VSH\[3\] analog/VOUTL analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[2\] analog/VOUTL analog/LSB_L_VSH\[3\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[2\] analog/VOUTL analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[2\] analog/LSB_L_VSH\[3\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[2\] analog/LSB_L_VSH\[3\] analog/VOUTL analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[2\] analog/VOUTL analog/LSB_L_VSH\[3\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[2\] analog/VOUTL analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[2\] analog/LSB_L_VSH\[3\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[2\] analog/LSB_L_VSH\[3\] analog/VOUTH analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[2\] analog/VOUTH analog/LSB_L_VSH\[3\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[2\] analog/VOUTH analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[2\] analog/LSB_L_VSH\[3\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[2\] analog/LSB_L_VSH\[3\] analog/VOUTH analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[2\] analog/VOUTH analog/LSB_L_VSH\[3\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[2\] analog/VOUTH analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[2\] analog/LSB_L_VSH\[3\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[2\] analog/LSB_L_VSH\[3\] analog/VOUTH analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[2\] analog/VOUTH analog/LSB_L_VSH\[3\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[2\] analog/VOUTH analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[2\] analog/LSB_L_VSH\[3\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[2\] analog/LSB_L_VSH\[3\] analog/VOUTH analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[2\] analog/VOUTH analog/LSB_L_VSH\[3\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[2\] analog/VOUTH analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[2\] analog/LSB_L_VSH\[3\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[0\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[10\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[11\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[12\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[13\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[14\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[15\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[16\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[17\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[18\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[19\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[1\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[20\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[21\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[22\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[23\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[2\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[3\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[4\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[5\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[6\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[7\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[8\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap\[9\].cap/impl
+ analog/LSB_L_VSH\[3\] analog/LSB_L_FL\[3\] analog/LSB_L_FL\[3\]
+ analog/LSB_L_FL\[3\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[3\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[3\] VREFL analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[3\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[3\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[3\] VREFL analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[3\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[3\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[3\] VREFL analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[3\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[3\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[3\] VREFL analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[3\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[3\] analog/LSB_L_VSH\[3\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1
+ analog/CRH\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2
+ analog/CRH\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1
+ analog/CRHB\[3\] analog/VOUTL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2
+ analog/CRHB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTL analog/VOUTL
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1
+ analog/CRL\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz2
+ analog/CRL\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1
+ analog/CRLB\[3\] analog/VOUTH analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2
+ analog/CRLB\[3\] analog/LSB_L_VSH\[4\] analog/VOUTH analog/VOUTH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[0\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[10\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[11\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[12\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[13\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[14\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[15\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[16\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[17\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[18\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[19\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[1\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[20\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[21\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[22\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[23\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[24\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[25\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[26\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[27\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[28\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[29\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[2\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[30\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[31\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[32\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[33\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[34\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[35\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[36\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[37\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[38\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[39\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[3\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[40\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[41\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[42\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[43\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[44\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[45\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[46\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[47\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[4\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[5\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[6\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[7\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[8\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap\[9\].cap/impl
+ analog/LSB_L_VSH\[4\] analog/LSB_L_FL\[4\] analog/LSB_L_FL\[4\]
+ analog/LSB_L_FL\[4\] AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[4\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[4\] VREFL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[4\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[4\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[4\] VREFL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[4\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[4\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[4\] VREFL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[4\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[4\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[4\] VREFL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[4\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[4\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[4\] VREFL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[4\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[4\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[4\] VREFL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[4\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[4\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[4\] VREFL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[4\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[4\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[4\] VREFL analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[4\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[4\] analog/LSB_L_VSH\[4\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/lsb_cdac_l.cdac_unit.CRH analog/LSB_L_VSH\[0\] analog/VOUTL
+ analog/LSB_L_VSH\[0\] AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/lsb_cdac_l.cdac_unit.CRH analog/VOUTL analog/LSB_L_VSH\[0\]
+ analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/lsb_cdac_l.cdac_unit.CRHB analog/VOUTL analog/LSB_L_VSH\[0\]
+ analog/LSB_L_VSH\[0\] AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/lsb_cdac_l.cdac_unit.CRHB analog/LSB_L_VSH\[0\] analog/VOUTL
+ analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/lsb_cdac_l.cdac_unit.CRH analog/LSB_L_VSH\[0\] analog/VOUTH
+ analog/LSB_L_VSH\[0\] AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/lsb_cdac_l.cdac_unit.CRH analog/VOUTH analog/LSB_L_VSH\[0\]
+ analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/lsb_cdac_l.cdac_unit.CRHB analog/VOUTH analog/LSB_L_VSH\[0\]
+ analog/LSB_L_VSH\[0\] AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/lsb_cdac_l.cdac_unit.CRHB analog/LSB_L_VSH\[0\] analog/VOUTH
+ analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.cap\[0\].cap/impl analog/LSB_L_VSH\[0\]
+ analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_unit.cap\[1\].cap/impl analog/LSB_L_VSH\[0\]
+ analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_unit.cap\[2\].cap/impl analog/LSB_L_VSH\[0\]
+ analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_unit.cap\[3\].cap/impl analog/LSB_L_VSH\[0\]
+ analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_unit.cap\[4\].cap/impl analog/LSB_L_VSH\[0\]
+ analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_unit.cap\[5\].cap/impl analog/LSB_L_VSH\[0\]
+ analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\] analog/LSB_L_FL\[0\]
+ AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CPRE VREFL analog/LSB_L_VSH\[0\] VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CPRE analog/LSB_L_VSH\[0\] VREFL analog/LSB_L_VSH\[0\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CPREB analog/LSB_L_VSH\[0\] VREFL VREFL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CPREB VREFL analog/LSB_L_VSH\[0\] analog/LSB_L_VSH\[0\]
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/lsb_cdac_l.tieh.impl AVDD VSS analog/lsb_cdac_l.cdac_unit.CRHB
+ sg13g2f_TIEH
Xanalog/lsb_cdac_l.tiel.impl AVDD VSS analog/lsb_cdac_l.cdac_unit.CRH
+ sg13g2f_TIEL
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_H_VSH VIP analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIP analog/MSB_H_VSH VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIP analog/MSB_H_VSH analog/MSB_H_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_H_VSH VIP VIP AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_h.cdac_unit.CRL analog/MSB_H_VSH VIN analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_h.cdac_unit.CRL VIN analog/MSB_H_VSH VIN AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_h.cdac_unit.CRLB VIN analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_h.cdac_unit.CRLB analog/MSB_H_VSH VIN VIN
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.cap\[0\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[10\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[11\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[12\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[13\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[14\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[15\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[16\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[17\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[18\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[19\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[1\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[20\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[21\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[22\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[23\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[24\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[25\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[26\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[27\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[28\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[29\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[2\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[30\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[31\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[32\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[33\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[34\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[35\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[36\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[37\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[38\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[39\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[3\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[40\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[41\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[42\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[43\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[44\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[45\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[46\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[47\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[48\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[49\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[4\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[50\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[51\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[52\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[53\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[54\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[55\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[56\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[57\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[58\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[59\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[5\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[60\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[61\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[62\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[63\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[64\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[65\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[66\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[67\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[68\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[69\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[6\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[70\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[71\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[72\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[73\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[74\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[75\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[76\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[77\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[78\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[79\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[7\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[80\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[81\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[82\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[83\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[84\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[85\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[86\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[87\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[88\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[89\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[8\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[90\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[91\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[92\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[93\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[94\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[95\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.cap\[9\].cap/impl analog/MSB_H_VSH
+ analog/MSB_H_FL analog/MSB_H_FL analog/MSB_H_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTH analog/MSB_H_VSH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_H_VSH analog/VOUTH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_H_VSH analog/VOUTH analog/VOUTH AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTH analog/MSB_H_VSH analog/MSB_H_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_h.tieh.impl AVDD VSS analog/msb_cdac_h.cdac_unit.CRLB
+ sg13g2f_TIEH
Xanalog/msb_cdac_h.tiel.impl AVDD VSS analog/msb_cdac_h.cdac_unit.CRL
+ sg13g2f_TIEL
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz1
+ analog/CPRE analog/MSB_L_VSH VIN analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2
+ analog/CPRE VIN analog/MSB_L_VSH VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz1
+ analog/CPREB VIN analog/MSB_L_VSH analog/MSB_L_VSH AVDD VSS
+ SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz2
+ analog/CPREB analog/MSB_L_VSH VIN VIN AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgn_lz1
+ analog/msb_cdac_l.cdac_unit.CRL analog/MSB_L_VSH VIP analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgn_lz2
+ analog/msb_cdac_l.cdac_unit.CRL VIP analog/MSB_L_VSH VIP AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz1
+ analog/msb_cdac_l.cdac_unit.CRLB VIP analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz2
+ analog/msb_cdac_l.cdac_unit.CRLB analog/MSB_L_VSH VIP VIP
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.cap\[0\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[10\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[11\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[12\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[13\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[14\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[15\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[16\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[17\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[18\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[19\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[1\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[20\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[21\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[22\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[23\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[24\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[25\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[26\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[27\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[28\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[29\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[2\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[30\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[31\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[32\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[33\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[34\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[35\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[36\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[37\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[38\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[39\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[3\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[40\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[41\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[42\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[43\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[44\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[45\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[46\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[47\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[48\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[49\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[4\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[50\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[51\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[52\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[53\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[54\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[55\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[56\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[57\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[58\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[59\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[5\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[60\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[61\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[62\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[63\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[64\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[65\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[66\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[67\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[68\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[69\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[6\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[70\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[71\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[72\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[73\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[74\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[75\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[76\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[77\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[78\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[79\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[7\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[80\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[81\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[82\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[83\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[84\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[85\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[86\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[87\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[88\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[89\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[8\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[90\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[91\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[92\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[93\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[94\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[95\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.cap\[9\].cap/impl analog/MSB_L_VSH
+ analog/MSB_L_FL analog/MSB_L_FL analog/MSB_L_FL AVDD VSS SARADC_CELL_INVX16_ASCAP
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz1
+ analog/CHOLD analog/VOUTL analog/MSB_L_VSH analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2
+ analog/CHOLD analog/MSB_L_VSH analog/VOUTL analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz1
+ analog/CHOLDB analog/MSB_L_VSH analog/VOUTL analog/VOUTL AVDD
+ VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz2
+ analog/CHOLDB analog/VOUTL analog/MSB_L_VSH analog/MSB_L_VSH
+ AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/msb_cdac_l.tieh.impl AVDD VSS analog/msb_cdac_l.cdac_unit.CRLB
+ sg13g2f_TIEH
Xanalog/msb_cdac_l.tiel.impl AVDD VSS analog/msb_cdac_l.cdac_unit.CRL
+ sg13g2f_TIEL
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz1 analog/CPRE
+ analog/VOUTH analog/VOUTL analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2 analog/CPRE
+ analog/VOUTL analog/VOUTH analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgp_lz1 analog/CPREB
+ analog/VOUTL analog/VOUTH analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgp_lz2 analog/CPREB
+ analog/VOUTH analog/VOUTL analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz1 analog/CPRE
+ analog/VOUTH analog/VOUTL analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2 analog/CPRE
+ analog/VOUTL analog/VOUTH analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgp_lz1 analog/CPREB
+ analog/VOUTL analog/VOUTH analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgp_lz2 analog/CPREB
+ analog/VOUTH analog/VOUTL analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgn_lz1 analog/CPRE
+ analog/VOUTH analog/VOUTL analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgn_lz2 analog/CPRE
+ analog/VOUTL analog/VOUTH analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgp_lz1 analog/CPREB
+ analog/VOUTL analog/VOUTH analog/VOUTH AVDD VSS SARADC_CELL_INVX0_ASSW
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgp_lz2 analog/CPREB
+ analog/VOUTH analog/VOUTL analog/VOUTL AVDD VSS SARADC_CELL_INVX0_ASSW
Xdigital/ins_051_ digital/state\[1\] digital/ins_017_ VSS
+ VDD sg13g2f_INVD1
Xdigital/ins_052_ digital/state\[0\] digital/ins_018_ VSS
+ VDD sg13g2f_INVD1
Xdigital/ins_053_ digital/mask\[0\] digital/ins_019_ VSS VDD
+ sg13g2f_INVD1
Xdigital/ins_054_ digital/mask\[1\] digital/ins_020_ VSS VDD
+ sg13g2f_INVD1
Xdigital/ins_055_ digital/mask\[2\] digital/ins_021_ VSS VDD
+ sg13g2f_INVD1
Xdigital/ins_056_ digital/mask\[3\] digital/ins_022_ VSS VDD
+ sg13g2f_INVD1
Xdigital/ins_057_ digital/mask\[4\] digital/ins_023_ VSS VDD
+ sg13g2f_INVD1
Xdigital/ins_058_ RST digital/ins_024_ VSS VDD sg13g2f_INVD1
Xdigital/ins_059_ RESULT[0] digital/ins_025_ VSS VDD sg13g2f_INVD1
Xdigital/ins_060_ RESULT[1] digital/ins_026_ VSS VDD sg13g2f_INVD1
Xdigital/ins_061_ RESULT[2] digital/ins_027_ VSS VDD sg13g2f_INVD1
Xdigital/ins_062_ RESULT[3] digital/ins_028_ VSS VDD sg13g2f_INVD1
Xdigital/ins_063_ RESULT[4] digital/ins_029_ VSS VDD sg13g2f_INVD1
Xdigital/ins_064_ digital/state\[1\] digital/ins_018_ RST
+ VDD VSS digital/ins_030_ sg13g2f_AOI21D1
Xdigital/ins_065_ digital/state\[1\] digital/ins_018_ RST
+ VDD VSS digital/ins_031_ sg13g2f_AO21D1
Xdigital/ins_066_ RST CMPO VDD VSS digital/ins_032_ sg13g2f_NR2D1
Xdigital/ins_067_ digital/mask\[0\] digital/ins_032_ RESULTN\[0\]
+ VDD VSS digital/ins_033_ sg13g2f_AO21D1
Xdigital/ins_068_ digital/ins_031_ digital/ins_033_ VDD VSS
+ digital/ins_000_ sg13g2f_AN2D1
Xdigital/ins_069_ digital/mask\[1\] digital/ins_032_ RESULTN\[1\]
+ VDD VSS digital/ins_034_ sg13g2f_AO21D1
Xdigital/ins_070_ digital/ins_031_ digital/ins_034_ VDD VSS
+ digital/ins_001_ sg13g2f_AN2D1
Xdigital/ins_071_ digital/mask\[2\] digital/ins_032_ RESULTN\[2\]
+ VDD VSS digital/ins_035_ sg13g2f_AO21D1
Xdigital/ins_072_ digital/ins_031_ digital/ins_035_ VDD VSS
+ digital/ins_002_ sg13g2f_AN2D1
Xdigital/ins_073_ digital/mask\[3\] digital/ins_032_ RESULTN\[3\]
+ VDD VSS digital/ins_036_ sg13g2f_AO21D1
Xdigital/ins_074_ digital/ins_031_ digital/ins_036_ VDD VSS
+ digital/ins_003_ sg13g2f_AN2D1
Xdigital/ins_075_ digital/mask\[4\] digital/ins_032_ RESULTN\[4\]
+ VDD VSS digital/ins_037_ sg13g2f_AO21D1
Xdigital/ins_076_ digital/ins_031_ digital/ins_037_ VDD VSS
+ digital/ins_004_ sg13g2f_AN2D1
Xdigital/ins_077_ digital/state\[1\] digital/ins_018_ digital/ins_024_
+ VDD VSS digital/ins_038_ sg13g2f_ND3D1
Xdigital/ins_078_ digital/ins_017_ digital/state\[0\] VDD
+ VSS SAMPLE sg13g2f_AN2D1
Xdigital/ins_079_ digital/ins_017_ digital/state\[0\] digital/ins_024_
+ VDD VSS digital/ins_039_ sg13g2f_ND3D1
Xdigital/ins_080_ digital/state\[1\] digital/state\[0\] VDD
+ VSS digital/ins_040_ sg13g2f_XNR2D1
Xdigital/ins_081_ RST digital/ins_040_ VDD VSS digital/ins_011_
+ sg13g2f_NR2D1
Xdigital/ins_082_ RST digital/ins_040_ digital/mask\[0\] VDD
+ VSS digital/ins_041_ sg13g2f_OAI21D1
Xdigital/ins_083_ digital/ins_020_ digital/ins_038_ digital/ins_041_
+ VDD VSS digital/ins_005_ sg13g2f_OAI21D1
Xdigital/ins_084_ RST digital/ins_040_ digital/mask\[1\] VDD
+ VSS digital/ins_042_ sg13g2f_OAI21D1
Xdigital/ins_085_ digital/ins_021_ digital/ins_038_ digital/ins_042_
+ VDD VSS digital/ins_006_ sg13g2f_OAI21D1
Xdigital/ins_086_ RST digital/ins_040_ digital/mask\[2\] VDD
+ VSS digital/ins_043_ sg13g2f_OAI21D1
Xdigital/ins_087_ digital/ins_022_ digital/ins_038_ digital/ins_043_
+ VDD VSS digital/ins_007_ sg13g2f_OAI21D1
Xdigital/ins_088_ RST digital/ins_040_ digital/mask\[3\] VDD
+ VSS digital/ins_044_ sg13g2f_OAI21D1
Xdigital/ins_089_ digital/ins_023_ digital/ins_038_ digital/ins_044_
+ VDD VSS digital/ins_008_ sg13g2f_OAI21D1
Xdigital/ins_090_ digital/ins_023_ digital/ins_011_ digital/ins_039_
+ VDD VSS digital/ins_009_ sg13g2f_OAI21D1
Xdigital/ins_091_ digital/ins_024_ GO digital/ins_040_ VDD
+ VSS digital/ins_045_ sg13g2f_ND3D1
Xdigital/ins_092_ digital/ins_019_ digital/ins_038_ digital/ins_045_
+ VDD VSS digital/ins_010_ sg13g2f_OAI21D1
Xdigital/ins_093_ digital/mask\[0\] digital/ins_024_ CMPO
+ VDD VSS digital/ins_046_ sg13g2f_ND3D1
Xdigital/ins_094_ digital/ins_025_ digital/ins_046_ digital/ins_030_
+ VDD VSS digital/ins_012_ sg13g2f_AOI21D1
Xdigital/ins_095_ digital/mask\[1\] digital/ins_024_ CMPO
+ VDD VSS digital/ins_047_ sg13g2f_ND3D1
Xdigital/ins_096_ digital/ins_026_ digital/ins_047_ digital/ins_030_
+ VDD VSS digital/ins_013_ sg13g2f_AOI21D1
Xdigital/ins_097_ digital/mask\[2\] digital/ins_024_ CMPO
+ VDD VSS digital/ins_048_ sg13g2f_ND3D1
Xdigital/ins_098_ digital/ins_027_ digital/ins_048_ digital/ins_030_
+ VDD VSS digital/ins_014_ sg13g2f_AOI21D1
Xdigital/ins_099_ digital/mask\[3\] digital/ins_024_ CMPO
+ VDD VSS digital/ins_049_ sg13g2f_ND3D1
Xdigital/ins_100_ digital/ins_028_ digital/ins_049_ digital/ins_030_
+ VDD VSS digital/ins_015_ sg13g2f_AOI21D1
Xdigital/ins_101_ digital/mask\[4\] digital/ins_024_ CMPO
+ VDD VSS digital/ins_050_ sg13g2f_ND3D1
Xdigital/ins_102_ digital/ins_029_ digital/ins_050_ digital/ins_030_
+ VDD VSS digital/ins_016_ sg13g2f_AOI21D1
Xdigital/ins_103_ digital/state\[1\] digital/state\[0\] VDD
+ VSS VALID sg13g2f_AN2D1
Xdigital/ins_104_ clknet_leaf_2_CLK digital/ins_000_ RESULTN\[0\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_105_ clknet_leaf_2_CLK digital/ins_001_ RESULTN\[1\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_106_ clknet_leaf_2_CLK digital/ins_002_ RESULTN\[2\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_107_ clknet_leaf_0_CLK digital/ins_003_ RESULTN\[3\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_108_ clknet_leaf_2_CLK digital/ins_004_ RESULTN\[4\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_109_ clknet_leaf_1_CLK digital/ins_005_ digital/mask\[0\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_110_ clknet_leaf_1_CLK digital/ins_006_ digital/mask\[1\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_111_ clknet_leaf_0_CLK digital/ins_007_ digital/mask\[2\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_112_ clknet_1_1__leaf_CLK digital/ins_008_ digital/mask\[3\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_113_ clknet_leaf_3_CLK digital/ins_009_ digital/mask\[4\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_114_ clknet_leaf_0_CLK digital/ins_010_ digital/state\[0\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_115_ clknet_leaf_0_CLK digital/ins_011_ digital/state\[1\]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_116_ clknet_leaf_3_CLK digital/ins_012_ RESULT[0]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_117_ clknet_leaf_1_CLK digital/ins_013_ RESULT[1]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_118_ clknet_leaf_1_CLK digital/ins_014_ RESULT[2]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_119_ clknet_leaf_3_CLK digital/ins_015_ RESULT[3]
+ VDD VSS sg13g2f_DFQD1
Xdigital/ins_120_ clknet_leaf_3_CLK digital/ins_016_ RESULT[4]
+ VDD VSS sg13g2f_DFQD1
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[0\].cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_unit_0_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_unit_0_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_unit_0_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_unit_0_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_unit_0_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_unit_0_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[1\].cdac_unit_1_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_1_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_2_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[2\].cdac_unit_3_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_1_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_2_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_3_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_4_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_5_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_6_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_h.cdac_bit\[3\].cdac_unit_7_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_0_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_0_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_0_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_0_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_0_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_0_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_1_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_1_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_1_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_1_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_1_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_1_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_2_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_2_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_2_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_2_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_2_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_2_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_3_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_3_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_3_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_3_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_3_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_3_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_4_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_4_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_4_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_4_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_4_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_4_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_5_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_5_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_5_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_5_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_5_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_5_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_6_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_6_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_6_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_6_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_6_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_6_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_7_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_7_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_7_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_7_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_7_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_7_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_8_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_8_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_8_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_8_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_8_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_8_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_9_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_9_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_9_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_9_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_9_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_9_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_10_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_10_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_10_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_10_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_10_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_10_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_11_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_11_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_11_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_11_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_11_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_11_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_12_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_12_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_12_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_12_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_12_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_12_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_13_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_13_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_13_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_13_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_13_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_13_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_14_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_14_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_14_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_14_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_14_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_14_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_15_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_15_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_15_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_15_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_h.cdac_unit_15_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_h.cdac_unit_15_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[0\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[1\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[2\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[3\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[4\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[5\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[6\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[7\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[8\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[9\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[10\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[11\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[12\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[13\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[14\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[15\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[16\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[17\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[18\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[19\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[20\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[21\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[22\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[23\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[24\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[25\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[26\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_h.dummy\[27\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgp_lz1_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgp_lz1_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz1_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz1_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgp_lz2_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgp_lz2_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[0\].impl/pgn_lz2_FILLA_7_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgp_lz1_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgp_lz1_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz1_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz1_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgp_lz2_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgp_lz2_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[1\].impl/pgn_lz2_FILLA_7_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgp_lz1_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgp_lz1_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgn_lz1_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgn_lz1_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgp_lz2_FILLM_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl.impl\[2\].impl/pgp_lz2_FILLM_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/sw_vouth2voutl_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLB_7_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPFILLA_7_0 SARADC_FILL1_NOPOWER
Xanalog/sw_vouth2voutl_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/sw_vouth2voutl_SW_TAPBB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/sw_vouth2voutl_SW_TAPAA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[0\].cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_unit_0_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_unit_0_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_unit_0_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_unit_0_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_unit_0_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_unit_0_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[1\].cdac_unit_1_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_1_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_2_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[2\].cdac_unit_3_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_1_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_2_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_3_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_4_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_5_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_6_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/lsb_cdac_l.cdac_bit\[3\].cdac_unit_7_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_0_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_0_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_0_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_0_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_0_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_0_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[1\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[1\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[1\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_1_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_1_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_1_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_1_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_1_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_1_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[2\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[2\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[2\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_2_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_2_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_2_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_2_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_2_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_2_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[3\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[3\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[3\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_3_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_3_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_3_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_3_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_3_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_3_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[4\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[4\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[4\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_4_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_4_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_4_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_4_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_4_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_4_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[5\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[5\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[5\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_5_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_5_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_5_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_5_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_5_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_5_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[6\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[6\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[6\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_6_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_6_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_6_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_6_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_6_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_6_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[7\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[7\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[7\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_7_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_7_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_7_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_7_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_7_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_7_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[8\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[8\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[8\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_8_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_8_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_8_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_8_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_8_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_8_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[9\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[9\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[9\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_9_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_9_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_9_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_9_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_9_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_9_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[10\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[10\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[10\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_10_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_10_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_10_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_10_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_10_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_10_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[11\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[11\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[11\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_11_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_11_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_11_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_11_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_11_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_11_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[12\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[12\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[12\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_12_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_12_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_12_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_12_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_12_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_12_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[13\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[13\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[13\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_13_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_13_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_13_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_13_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_13_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_13_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[14\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[14\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[14\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_14_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_14_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_14_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_14_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_14_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_14_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.vi2cap\[15\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2vouth\[15\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit.cap2voutl\[15\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_CAP_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_15_CAP_TAPB_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_15_CAP_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_CAP_TAPFILLB_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_CAP_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_CAP_TAPFILLA_0_1 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_CAP_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_15_CAP_TAPA_0_1 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_15_SW_TAPB_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/msb_cdac_l.cdac_unit_15_SW_TAPFILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_SW_TAPFILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/msb_cdac_l.cdac_unit_15_SW_TAPA_0_0 AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[0\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[1\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[2\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[3\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[4\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[5\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[6\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[7\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[8\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_SW_TAPB_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[9\].dummy.cdac_unit_0_SW_TAPA_0_0 AVDD
+ VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[10\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[11\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[12\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[13\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[14\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[15\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[16\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[17\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_CAP_TAPAA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[18\].dummy.cdac_unit_0_SW_TAPAA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[19\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[20\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[21\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[22\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[23\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[24\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[25\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[26\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.vi2cap\[0\].sw_vi2cap/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_2_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_3_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_4_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_5_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_6_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2vouth\[0\].sw_cap2vouth/pgn_lz2_FILLA_7_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgn_lz1_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit.cap2voutl\[0\].sw_cap2voutl/pgp_lz2_FILLM_1_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLB_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLB_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLB_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLB_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLB_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLB_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLB_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLA_0_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLA_1_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLA_2_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLA_3_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLA_4_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLA_5_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_FILLA_6_0 SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPFILLB_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPFILLA_0_1
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPA_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_SW_TAPB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_SW_TAPFILLB_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_SW_TAPFILLA_0_0
+ SARADC_FILL1_NOPOWER
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_SW_TAPA_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_CAP_TAPBB_0_1
+ AVDD VSS SARADC_FILLTIE2
Xanalog/dummy_l.dummy\[27\].dummy.cdac_unit_0_SW_TAPBB_0_0
+ AVDD VSS SARADC_FILLTIE2
Xtapcell_up_inst_1 AVDD VSS sg13g2f_TAPCELL
Xtapcell_dw_inst_1 AVDD VSS sg13g2f_TAPCELL
Xtapcell_up_inst_3 AVDD VSS sg13g2f_TAPCELL
Xtapcell_dw_inst_3 AVDD VSS sg13g2f_TAPCELL
Xtapcell_up_inst_7 AVDD VSS sg13g2f_TAPCELL
Xtapcell_dw_inst_7 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_25_ANALOG_2_Left_0 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_26_ANALOG_2_Left_1 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_27_ANALOG_2_Left_2 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_22_ANALOG_Left_3 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_23_ANALOG_Left_4 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_24_ANALOG_Left_5 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_25_ANALOG_2_Right_6 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_22_ANALOG_Right_7 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_23_ANALOG_Right_8 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_24_ANALOG_Right_9 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_26_ANALOG_2_Right_10 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_27_ANALOG_2_Right_11 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_28_ANALOG_Right_12 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_29_ANALOG_Right_13 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_30_ANALOG_Right_14 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_28_ANALOG_Left_15 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_29_ANALOG_Left_16 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_30_ANALOG_Left_17 AVDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_52_2_Right_18 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_51_2_Right_19 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_50_2_Right_20 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_49_2_Right_21 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_48_2_Right_22 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_47_2_Right_23 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_46_2_Right_24 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_45_2_Right_25 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_44_2_Right_26 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_43_2_Right_27 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_42_2_Right_28 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_41_2_Right_29 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_40_2_Right_30 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_39_2_Right_31 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_38_2_Right_32 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_37_2_Right_33 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_36_2_Right_34 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_35_2_Right_35 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_34_2_Right_36 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_33_2_Right_37 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_32_2_Right_38 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_31_2_Right_39 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_30_2_Right_40 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_29_2_Right_41 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_28_2_Right_42 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_27_2_Right_43 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_26_2_Right_44 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_25_2_Right_45 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_24_2_Right_46 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_23_2_Right_47 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_22_2_Right_48 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_21_2_Right_49 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_20_2_Right_50 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_19_2_Right_51 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_18_2_Right_52 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_17_2_Right_53 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_16_2_Right_54 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_15_2_Right_55 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_14_2_Right_56 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_13_2_Right_57 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_12_2_Right_58 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_11_2_Right_59 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_10_2_Right_60 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_9_2_Right_61 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_8_2_Right_62 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_7_2_Right_63 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_6_2_Right_64 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_5_2_Right_65 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_4_2_Right_66 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_3_2_Right_67 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_2_2_Right_68 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_1_2_Right_69 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_0_2_Right_70 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_52_2_Left_71 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_51_2_Left_72 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_50_2_Left_73 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_49_2_Left_74 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_48_2_Left_75 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_47_2_Left_76 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_46_2_Left_77 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_45_2_Left_78 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_44_2_Left_79 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_43_2_Left_80 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_42_2_Left_81 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_41_2_Left_82 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_40_2_Left_83 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_39_2_Left_84 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_38_2_Left_85 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_37_2_Left_86 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_36_2_Left_87 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_35_2_Left_88 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_34_2_Left_89 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_33_2_Left_90 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_32_2_Left_91 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_31_2_Left_92 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_30_2_Left_93 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_29_2_Left_94 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_28_2_Left_95 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_27_2_Left_96 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_26_2_Left_97 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_25_2_Left_98 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_24_2_Left_99 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_23_2_Left_100 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_22_2_Left_101 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_21_2_Left_102 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_20_2_Left_103 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_19_2_Left_104 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_18_2_Left_105 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_17_2_Left_106 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_16_2_Left_107 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_15_2_Left_108 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_14_2_Left_109 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_13_2_Left_110 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_12_2_Left_111 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_11_2_Left_112 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_10_2_Left_113 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_9_2_Left_114 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_8_2_Left_115 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_7_2_Left_116 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_6_2_Left_117 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_5_2_Left_118 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_4_2_Left_119 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_3_2_Left_120 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_2_2_Left_121 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_1_2_Left_122 VDD VSS sg13g2f_TAPCELL
XPHY_EDGE_ROW_0_2_Left_123 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_25_ANALOG_2_124 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_25_ANALOG_2_125 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_25_ANALOG_2_126 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_25_ANALOG_2_127 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_128 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_129 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_130 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_131 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_132 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_133 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_134 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_135 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_136 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_137 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_ANALOG_138 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_23_ANALOG_139 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_23_ANALOG_140 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_23_ANALOG_141 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_23_ANALOG_142 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_23_ANALOG_143 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_144 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_145 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_146 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_147 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_148 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_149 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_150 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_151 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_152 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_153 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_ANALOG_154 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_26_ANALOG_2_155 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_26_ANALOG_2_156 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_26_ANALOG_2_157 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_26_ANALOG_2_158 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_27_ANALOG_2_159 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_27_ANALOG_2_160 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_27_ANALOG_2_161 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_162 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_163 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_164 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_165 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_166 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_167 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_168 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_169 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_170 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_171 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_ANALOG_172 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_29_ANALOG_173 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_29_ANALOG_174 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_29_ANALOG_175 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_29_ANALOG_176 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_29_ANALOG_177 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_178 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_179 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_180 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_181 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_182 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_183 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_184 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_185 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_186 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_187 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_ANALOG_188 AVDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_52_2_189 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_50_2_190 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_48_2_191 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_46_2_192 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_44_2_193 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_42_2_194 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_40_2_195 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_38_2_196 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_36_2_197 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_34_2_198 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_32_2_199 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_30_2_200 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_28_2_201 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_26_2_202 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_24_2_203 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_22_2_204 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_20_2_205 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_18_2_206 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_16_2_207 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_14_2_208 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_12_2_209 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_10_2_210 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_8_2_211 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_6_2_212 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_4_2_213 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_2_2_214 VDD VSS sg13g2f_TAPCELL
XTAP_TAPCELL_ROW_0_2_215 VDD VSS sg13g2f_TAPCELL
Xclkbuf_regs_0_CLK CLK VDD VSS CLK_regs sg13g2f_BUFFD1
Xclkbuf_leaf_0_CLK clknet_1_1__leaf_CLK VDD VSS clknet_leaf_0_CLK
+ sg13g2f_BUFFD1
Xclkbuf_leaf_1_CLK clknet_1_1__leaf_CLK VDD VSS clknet_leaf_1_CLK
+ sg13g2f_BUFFD1
Xclkbuf_leaf_2_CLK clknet_1_0__leaf_CLK VDD VSS clknet_leaf_2_CLK
+ sg13g2f_BUFFD1
Xclkbuf_leaf_3_CLK clknet_1_0__leaf_CLK VDD VSS clknet_leaf_3_CLK
+ sg13g2f_BUFFD1
Xclkbuf_0_CLK CLK VDD VSS clknet_0_CLK sg13g2f_BUFFD1
Xclkbuf_1_0__f_CLK clknet_0_CLK VDD VSS clknet_1_0__leaf_CLK
+ sg13g2f_BUFFD1
Xclkbuf_1_1__f_CLK clknet_0_CLK VDD VSS clknet_1_1__leaf_CLK
+ sg13g2f_BUFFD1
Xclkload0 clknet_1_0__leaf_CLK _unconnected_0 VSS VDD sg13g2f_INVD1
Xclkbuf_0_CLK_regs CLK_regs VDD VSS clknet_0_CLK_regs sg13g2f_BUFFD1
Xclkbuf_1_0__f_CLK_regs clknet_0_CLK_regs VDD VSS clknet_1_0__leaf_CLK_regs
+ sg13g2f_BUFFD1
XFILLER_0_1390 VDD VSS sg13g2f_FILL8
XFILLER_0_1398 VDD VSS sg13g2f_FILL8
XFILLER_0_1406 VDD VSS sg13g2f_FILL8
XFILLER_0_1414 VDD VSS sg13g2f_FILL8
XFILLER_0_1422 VDD VSS sg13g2f_FILL8
XFILLER_0_1430 VDD VSS sg13g2f_FILL8
XFILLER_0_1438 VDD VSS sg13g2f_FILL8
XFILLER_0_1446 VDD VSS sg13g2f_FILL8
XFILLER_0_1454 VDD VSS sg13g2f_FILL8
XFILLER_0_1462 VDD VSS sg13g2f_FILL8
XFILLER_0_1470 VDD VSS sg13g2f_FILL8
XFILLER_0_1478 VDD VSS sg13g2f_FILL8
XFILLER_0_1486 VDD VSS sg13g2f_FILL8
XFILLER_0_1494 VDD VSS sg13g2f_FILL1
XFILLER_0_1502 VDD VSS sg13g2f_FILL8
XFILLER_0_1510 VDD VSS sg13g2f_FILL8
XFILLER_0_1518 VDD VSS sg13g2f_FILL8
XFILLER_0_1526 VDD VSS sg13g2f_FILL8
XFILLER_0_1534 VDD VSS sg13g2f_FILL8
XFILLER_0_1542 VDD VSS sg13g2f_FILL8
XFILLER_0_1550 VDD VSS sg13g2f_FILL1
XFILLER_1_1390 VDD VSS sg13g2f_FILL8
XFILLER_1_1398 VDD VSS sg13g2f_FILL8
XFILLER_1_1406 VDD VSS sg13g2f_FILL8
XFILLER_1_1414 VDD VSS sg13g2f_FILL8
XFILLER_1_1422 VDD VSS sg13g2f_FILL8
XFILLER_1_1430 VDD VSS sg13g2f_FILL8
XFILLER_1_1438 VDD VSS sg13g2f_FILL8
XFILLER_1_1446 VDD VSS sg13g2f_FILL8
XFILLER_1_1454 VDD VSS sg13g2f_FILL8
XFILLER_1_1462 VDD VSS sg13g2f_FILL8
XFILLER_1_1470 VDD VSS sg13g2f_FILL8
XFILLER_1_1478 VDD VSS sg13g2f_FILL8
XFILLER_1_1486 VDD VSS sg13g2f_FILL8
XFILLER_1_1494 VDD VSS sg13g2f_FILL8
XFILLER_1_1502 VDD VSS sg13g2f_FILL8
XFILLER_1_1510 VDD VSS sg13g2f_FILL4
XFILLER_1_1514 VDD VSS sg13g2f_FILL1
XFILLER_1_1526 VDD VSS sg13g2f_FILL8
XFILLER_1_1534 VDD VSS sg13g2f_FILL8
XFILLER_1_1542 VDD VSS sg13g2f_FILL8
XFILLER_1_1550 VDD VSS sg13g2f_FILL1
XFILLER_2_1390 VDD VSS sg13g2f_FILL8
XFILLER_2_1398 VDD VSS sg13g2f_FILL8
XFILLER_2_1406 VDD VSS sg13g2f_FILL8
XFILLER_2_1414 VDD VSS sg13g2f_FILL8
XFILLER_2_1422 VDD VSS sg13g2f_FILL8
XFILLER_2_1430 VDD VSS sg13g2f_FILL8
XFILLER_2_1438 VDD VSS sg13g2f_FILL8
XFILLER_2_1446 VDD VSS sg13g2f_FILL8
XFILLER_2_1454 VDD VSS sg13g2f_FILL8
XFILLER_2_1462 VDD VSS sg13g2f_FILL8
XFILLER_2_1470 VDD VSS sg13g2f_FILL8
XFILLER_2_1478 VDD VSS sg13g2f_FILL8
XFILLER_2_1486 VDD VSS sg13g2f_FILL8
XFILLER_2_1494 VDD VSS sg13g2f_FILL4
XFILLER_2_1505 VDD VSS sg13g2f_FILL8
XFILLER_2_1513 VDD VSS sg13g2f_FILL8
XFILLER_2_1521 VDD VSS sg13g2f_FILL8
XFILLER_2_1529 VDD VSS sg13g2f_FILL8
XFILLER_2_1537 VDD VSS sg13g2f_FILL8
XFILLER_2_1545 VDD VSS sg13g2f_FILL4
XFILLER_2_1549 VDD VSS sg13g2f_FILL2
XFILLER_3_1390 VDD VSS sg13g2f_FILL8
XFILLER_3_1398 VDD VSS sg13g2f_FILL8
XFILLER_3_1406 VDD VSS sg13g2f_FILL8
XFILLER_3_1414 VDD VSS sg13g2f_FILL8
XFILLER_3_1422 VDD VSS sg13g2f_FILL8
XFILLER_3_1430 VDD VSS sg13g2f_FILL8
XFILLER_3_1438 VDD VSS sg13g2f_FILL8
XFILLER_3_1446 VDD VSS sg13g2f_FILL8
XFILLER_3_1454 VDD VSS sg13g2f_FILL8
XFILLER_3_1462 VDD VSS sg13g2f_FILL8
XFILLER_3_1470 VDD VSS sg13g2f_FILL8
XFILLER_3_1478 VDD VSS sg13g2f_FILL8
XFILLER_3_1486 VDD VSS sg13g2f_FILL8
XFILLER_3_1494 VDD VSS sg13g2f_FILL8
XFILLER_3_1502 VDD VSS sg13g2f_FILL2
XFILLER_3_1504 VDD VSS sg13g2f_FILL1
XFILLER_3_1537 VDD VSS sg13g2f_FILL8
XFILLER_3_1545 VDD VSS sg13g2f_FILL4
XFILLER_3_1549 VDD VSS sg13g2f_FILL2
XFILLER_4_1390 VDD VSS sg13g2f_FILL8
XFILLER_4_1398 VDD VSS sg13g2f_FILL8
XFILLER_4_1406 VDD VSS sg13g2f_FILL8
XFILLER_4_1414 VDD VSS sg13g2f_FILL8
XFILLER_4_1422 VDD VSS sg13g2f_FILL8
XFILLER_4_1430 VDD VSS sg13g2f_FILL8
XFILLER_4_1438 VDD VSS sg13g2f_FILL8
XFILLER_4_1446 VDD VSS sg13g2f_FILL8
XFILLER_4_1454 VDD VSS sg13g2f_FILL8
XFILLER_4_1462 VDD VSS sg13g2f_FILL8
XFILLER_4_1470 VDD VSS sg13g2f_FILL8
XFILLER_4_1478 VDD VSS sg13g2f_FILL8
XFILLER_4_1486 VDD VSS sg13g2f_FILL8
XFILLER_4_1494 VDD VSS sg13g2f_FILL4
XFILLER_4_1505 VDD VSS sg13g2f_FILL8
XFILLER_4_1513 VDD VSS sg13g2f_FILL2
XFILLER_4_1515 VDD VSS sg13g2f_FILL1
XFILLER_4_1527 VDD VSS sg13g2f_FILL8
XFILLER_4_1535 VDD VSS sg13g2f_FILL8
XFILLER_4_1543 VDD VSS sg13g2f_FILL8
XFILLER_5_1390 VDD VSS sg13g2f_FILL8
XFILLER_5_1398 VDD VSS sg13g2f_FILL8
XFILLER_5_1406 VDD VSS sg13g2f_FILL8
XFILLER_5_1414 VDD VSS sg13g2f_FILL8
XFILLER_5_1422 VDD VSS sg13g2f_FILL8
XFILLER_5_1430 VDD VSS sg13g2f_FILL8
XFILLER_5_1438 VDD VSS sg13g2f_FILL8
XFILLER_5_1446 VDD VSS sg13g2f_FILL8
XFILLER_5_1454 VDD VSS sg13g2f_FILL8
XFILLER_5_1462 VDD VSS sg13g2f_FILL8
XFILLER_5_1470 VDD VSS sg13g2f_FILL8
XFILLER_5_1478 VDD VSS sg13g2f_FILL8
XFILLER_5_1486 VDD VSS sg13g2f_FILL8
XFILLER_5_1494 VDD VSS sg13g2f_FILL4
XFILLER_5_1498 VDD VSS sg13g2f_FILL2
XFILLER_5_1500 VDD VSS sg13g2f_FILL1
XFILLER_5_1543 VDD VSS sg13g2f_FILL8
XFILLER_6_1390 VDD VSS sg13g2f_FILL8
XFILLER_6_1398 VDD VSS sg13g2f_FILL8
XFILLER_6_1406 VDD VSS sg13g2f_FILL8
XFILLER_6_1414 VDD VSS sg13g2f_FILL8
XFILLER_6_1422 VDD VSS sg13g2f_FILL8
XFILLER_6_1430 VDD VSS sg13g2f_FILL8
XFILLER_6_1438 VDD VSS sg13g2f_FILL8
XFILLER_6_1446 VDD VSS sg13g2f_FILL8
XFILLER_6_1454 VDD VSS sg13g2f_FILL8
XFILLER_6_1462 VDD VSS sg13g2f_FILL8
XFILLER_6_1470 VDD VSS sg13g2f_FILL8
XFILLER_6_1478 VDD VSS sg13g2f_FILL8
XFILLER_6_1486 VDD VSS sg13g2f_FILL8
XFILLER_6_1494 VDD VSS sg13g2f_FILL4
XFILLER_6_1547 VDD VSS sg13g2f_FILL4
XFILLER_7_1390 VDD VSS sg13g2f_FILL8
XFILLER_7_1398 VDD VSS sg13g2f_FILL8
XFILLER_7_1406 VDD VSS sg13g2f_FILL8
XFILLER_7_1414 VDD VSS sg13g2f_FILL8
XFILLER_7_1422 VDD VSS sg13g2f_FILL8
XFILLER_7_1430 VDD VSS sg13g2f_FILL8
XFILLER_7_1438 VDD VSS sg13g2f_FILL8
XFILLER_7_1446 VDD VSS sg13g2f_FILL8
XFILLER_7_1454 VDD VSS sg13g2f_FILL8
XFILLER_7_1462 VDD VSS sg13g2f_FILL8
XFILLER_7_1470 VDD VSS sg13g2f_FILL8
XFILLER_7_1478 VDD VSS sg13g2f_FILL8
XFILLER_7_1486 VDD VSS sg13g2f_FILL8
XFILLER_7_1494 VDD VSS sg13g2f_FILL8
XFILLER_7_1502 VDD VSS sg13g2f_FILL8
XFILLER_7_1510 VDD VSS sg13g2f_FILL8
XFILLER_7_1518 VDD VSS sg13g2f_FILL8
XFILLER_7_1526 VDD VSS sg13g2f_FILL8
XFILLER_7_1534 VDD VSS sg13g2f_FILL8
XFILLER_7_1542 VDD VSS sg13g2f_FILL8
XFILLER_7_1550 VDD VSS sg13g2f_FILL1
XFILLER_8_1390 VDD VSS sg13g2f_FILL8
XFILLER_8_1398 VDD VSS sg13g2f_FILL8
XFILLER_8_1406 VDD VSS sg13g2f_FILL8
XFILLER_8_1414 VDD VSS sg13g2f_FILL8
XFILLER_8_1422 VDD VSS sg13g2f_FILL8
XFILLER_8_1430 VDD VSS sg13g2f_FILL8
XFILLER_8_1438 VDD VSS sg13g2f_FILL8
XFILLER_8_1446 VDD VSS sg13g2f_FILL8
XFILLER_8_1454 VDD VSS sg13g2f_FILL8
XFILLER_8_1462 VDD VSS sg13g2f_FILL8
XFILLER_8_1470 VDD VSS sg13g2f_FILL8
XFILLER_8_1478 VDD VSS sg13g2f_FILL8
XFILLER_8_1486 VDD VSS sg13g2f_FILL8
XFILLER_8_1494 VDD VSS sg13g2f_FILL4
XFILLER_8_1547 VDD VSS sg13g2f_FILL4
XFILLER_9_1390 VDD VSS sg13g2f_FILL8
XFILLER_9_1398 VDD VSS sg13g2f_FILL8
XFILLER_9_1406 VDD VSS sg13g2f_FILL8
XFILLER_9_1414 VDD VSS sg13g2f_FILL8
XFILLER_9_1422 VDD VSS sg13g2f_FILL8
XFILLER_9_1430 VDD VSS sg13g2f_FILL8
XFILLER_9_1438 VDD VSS sg13g2f_FILL8
XFILLER_9_1446 VDD VSS sg13g2f_FILL8
XFILLER_9_1454 VDD VSS sg13g2f_FILL8
XFILLER_9_1462 VDD VSS sg13g2f_FILL8
XFILLER_9_1470 VDD VSS sg13g2f_FILL8
XFILLER_9_1478 VDD VSS sg13g2f_FILL8
XFILLER_9_1486 VDD VSS sg13g2f_FILL8
XFILLER_9_1494 VDD VSS sg13g2f_FILL8
XFILLER_9_1502 VDD VSS sg13g2f_FILL8
XFILLER_9_1510 VDD VSS sg13g2f_FILL8
XFILLER_9_1518 VDD VSS sg13g2f_FILL8
XFILLER_9_1526 VDD VSS sg13g2f_FILL8
XFILLER_9_1534 VDD VSS sg13g2f_FILL8
XFILLER_9_1542 VDD VSS sg13g2f_FILL8
XFILLER_9_1550 VDD VSS sg13g2f_FILL1
XFILLER_10_1390 VDD VSS sg13g2f_FILL8
XFILLER_10_1398 VDD VSS sg13g2f_FILL8
XFILLER_10_1406 VDD VSS sg13g2f_FILL8
XFILLER_10_1414 VDD VSS sg13g2f_FILL8
XFILLER_10_1422 VDD VSS sg13g2f_FILL8
XFILLER_10_1430 VDD VSS sg13g2f_FILL8
XFILLER_10_1438 VDD VSS sg13g2f_FILL8
XFILLER_10_1446 VDD VSS sg13g2f_FILL8
XFILLER_10_1454 VDD VSS sg13g2f_FILL8
XFILLER_10_1462 VDD VSS sg13g2f_FILL8
XFILLER_10_1470 VDD VSS sg13g2f_FILL8
XFILLER_10_1478 VDD VSS sg13g2f_FILL8
XFILLER_10_1486 VDD VSS sg13g2f_FILL8
XFILLER_10_1494 VDD VSS sg13g2f_FILL4
XFILLER_10_1538 VDD VSS sg13g2f_FILL8
XFILLER_10_1546 VDD VSS sg13g2f_FILL4
XFILLER_10_1550 VDD VSS sg13g2f_FILL1
XFILLER_11_1390 VDD VSS sg13g2f_FILL8
XFILLER_11_1398 VDD VSS sg13g2f_FILL8
XFILLER_11_1406 VDD VSS sg13g2f_FILL8
XFILLER_11_1414 VDD VSS sg13g2f_FILL8
XFILLER_11_1422 VDD VSS sg13g2f_FILL8
XFILLER_11_1430 VDD VSS sg13g2f_FILL8
XFILLER_11_1438 VDD VSS sg13g2f_FILL8
XFILLER_11_1446 VDD VSS sg13g2f_FILL8
XFILLER_11_1454 VDD VSS sg13g2f_FILL8
XFILLER_11_1462 VDD VSS sg13g2f_FILL8
XFILLER_11_1470 VDD VSS sg13g2f_FILL8
XFILLER_11_1478 VDD VSS sg13g2f_FILL4
XFILLER_11_1482 VDD VSS sg13g2f_FILL2
XFILLER_11_1484 VDD VSS sg13g2f_FILL1
XFILLER_11_1548 VDD VSS sg13g2f_FILL2
XFILLER_11_1550 VDD VSS sg13g2f_FILL1
XFILLER_12_1390 VDD VSS sg13g2f_FILL8
XFILLER_12_1398 VDD VSS sg13g2f_FILL8
XFILLER_12_1406 VDD VSS sg13g2f_FILL8
XFILLER_12_1414 VDD VSS sg13g2f_FILL8
XFILLER_12_1422 VDD VSS sg13g2f_FILL8
XFILLER_12_1430 VDD VSS sg13g2f_FILL8
XFILLER_12_1438 VDD VSS sg13g2f_FILL8
XFILLER_12_1446 VDD VSS sg13g2f_FILL8
XFILLER_12_1454 VDD VSS sg13g2f_FILL8
XFILLER_12_1462 VDD VSS sg13g2f_FILL8
XFILLER_12_1470 VDD VSS sg13g2f_FILL8
XFILLER_12_1478 VDD VSS sg13g2f_FILL8
XFILLER_12_1486 VDD VSS sg13g2f_FILL8
XFILLER_12_1494 VDD VSS sg13g2f_FILL4
XFILLER_12_1505 VDD VSS sg13g2f_FILL4
XFILLER_12_1536 VDD VSS sg13g2f_FILL2
XFILLER_12_1538 VDD VSS sg13g2f_FILL1
XFILLER_12_1547 VDD VSS sg13g2f_FILL4
XFILLER_13_1390 VDD VSS sg13g2f_FILL8
XFILLER_13_1398 VDD VSS sg13g2f_FILL8
XFILLER_13_1406 VDD VSS sg13g2f_FILL8
XFILLER_13_1414 VDD VSS sg13g2f_FILL8
XFILLER_13_1422 VDD VSS sg13g2f_FILL8
XFILLER_13_1430 VDD VSS sg13g2f_FILL8
XFILLER_13_1438 VDD VSS sg13g2f_FILL8
XFILLER_13_1446 VDD VSS sg13g2f_FILL8
XFILLER_13_1454 VDD VSS sg13g2f_FILL8
XFILLER_13_1462 VDD VSS sg13g2f_FILL8
XFILLER_13_1470 VDD VSS sg13g2f_FILL8
XFILLER_13_1478 VDD VSS sg13g2f_FILL8
XFILLER_13_1486 VDD VSS sg13g2f_FILL8
XFILLER_13_1494 VDD VSS sg13g2f_FILL4
XFILLER_13_1498 VDD VSS sg13g2f_FILL2
XFILLER_13_1542 VDD VSS sg13g2f_FILL8
XFILLER_13_1550 VDD VSS sg13g2f_FILL1
XFILLER_14_1390 VDD VSS sg13g2f_FILL8
XFILLER_14_1398 VDD VSS sg13g2f_FILL8
XFILLER_14_1406 VDD VSS sg13g2f_FILL8
XFILLER_14_1414 VDD VSS sg13g2f_FILL8
XFILLER_14_1422 VDD VSS sg13g2f_FILL8
XFILLER_14_1430 VDD VSS sg13g2f_FILL8
XFILLER_14_1438 VDD VSS sg13g2f_FILL8
XFILLER_14_1446 VDD VSS sg13g2f_FILL8
XFILLER_14_1454 VDD VSS sg13g2f_FILL8
XFILLER_14_1462 VDD VSS sg13g2f_FILL8
XFILLER_14_1470 VDD VSS sg13g2f_FILL8
XFILLER_14_1478 VDD VSS sg13g2f_FILL4
XFILLER_14_1482 VDD VSS sg13g2f_FILL2
XFILLER_14_1484 VDD VSS sg13g2f_FILL1
XFILLER_14_1547 VDD VSS sg13g2f_FILL4
XFILLER_15_1390 VDD VSS sg13g2f_FILL8
XFILLER_15_1398 VDD VSS sg13g2f_FILL8
XFILLER_15_1406 VDD VSS sg13g2f_FILL8
XFILLER_15_1414 VDD VSS sg13g2f_FILL8
XFILLER_15_1422 VDD VSS sg13g2f_FILL8
XFILLER_15_1430 VDD VSS sg13g2f_FILL8
XFILLER_15_1438 VDD VSS sg13g2f_FILL8
XFILLER_15_1446 VDD VSS sg13g2f_FILL8
XFILLER_15_1454 VDD VSS sg13g2f_FILL8
XFILLER_15_1462 VDD VSS sg13g2f_FILL8
XFILLER_15_1470 VDD VSS sg13g2f_FILL8
XFILLER_15_1478 VDD VSS sg13g2f_FILL8
XFILLER_15_1486 VDD VSS sg13g2f_FILL8
XFILLER_15_1494 VDD VSS sg13g2f_FILL8
XFILLER_15_1502 VDD VSS sg13g2f_FILL8
XFILLER_15_1510 VDD VSS sg13g2f_FILL4
XFILLER_15_1525 VDD VSS sg13g2f_FILL8
XFILLER_15_1533 VDD VSS sg13g2f_FILL8
XFILLER_15_1541 VDD VSS sg13g2f_FILL8
XFILLER_15_1549 VDD VSS sg13g2f_FILL2
XFILLER_16_1390 VDD VSS sg13g2f_FILL8
XFILLER_16_1398 VDD VSS sg13g2f_FILL8
XFILLER_16_1406 VDD VSS sg13g2f_FILL8
XFILLER_16_1414 VDD VSS sg13g2f_FILL8
XFILLER_16_1422 VDD VSS sg13g2f_FILL8
XFILLER_16_1430 VDD VSS sg13g2f_FILL8
XFILLER_16_1438 VDD VSS sg13g2f_FILL8
XFILLER_16_1446 VDD VSS sg13g2f_FILL8
XFILLER_16_1454 VDD VSS sg13g2f_FILL8
XFILLER_16_1462 VDD VSS sg13g2f_FILL8
XFILLER_16_1470 VDD VSS sg13g2f_FILL8
XFILLER_16_1478 VDD VSS sg13g2f_FILL8
XFILLER_16_1486 VDD VSS sg13g2f_FILL8
XFILLER_16_1494 VDD VSS sg13g2f_FILL4
XFILLER_16_1547 VDD VSS sg13g2f_FILL4
XFILLER_17_1390 VDD VSS sg13g2f_FILL8
XFILLER_17_1398 VDD VSS sg13g2f_FILL8
XFILLER_17_1406 VDD VSS sg13g2f_FILL8
XFILLER_17_1414 VDD VSS sg13g2f_FILL8
XFILLER_17_1422 VDD VSS sg13g2f_FILL8
XFILLER_17_1430 VDD VSS sg13g2f_FILL8
XFILLER_17_1438 VDD VSS sg13g2f_FILL8
XFILLER_17_1446 VDD VSS sg13g2f_FILL8
XFILLER_17_1454 VDD VSS sg13g2f_FILL8
XFILLER_17_1462 VDD VSS sg13g2f_FILL8
XFILLER_17_1470 VDD VSS sg13g2f_FILL8
XFILLER_17_1478 VDD VSS sg13g2f_FILL8
XFILLER_17_1486 VDD VSS sg13g2f_FILL8
XFILLER_17_1494 VDD VSS sg13g2f_FILL8
XFILLER_17_1502 VDD VSS sg13g2f_FILL8
XFILLER_17_1510 VDD VSS sg13g2f_FILL8
XFILLER_17_1518 VDD VSS sg13g2f_FILL8
XFILLER_17_1526 VDD VSS sg13g2f_FILL8
XFILLER_17_1534 VDD VSS sg13g2f_FILL8
XFILLER_17_1542 VDD VSS sg13g2f_FILL8
XFILLER_17_1550 VDD VSS sg13g2f_FILL1
XFILLER_18_1390 VDD VSS sg13g2f_FILL8
XFILLER_18_1398 VDD VSS sg13g2f_FILL8
XFILLER_18_1406 VDD VSS sg13g2f_FILL8
XFILLER_18_1414 VDD VSS sg13g2f_FILL8
XFILLER_18_1422 VDD VSS sg13g2f_FILL8
XFILLER_18_1430 VDD VSS sg13g2f_FILL8
XFILLER_18_1438 VDD VSS sg13g2f_FILL8
XFILLER_18_1446 VDD VSS sg13g2f_FILL8
XFILLER_18_1454 VDD VSS sg13g2f_FILL8
XFILLER_18_1462 VDD VSS sg13g2f_FILL8
XFILLER_18_1470 VDD VSS sg13g2f_FILL8
XFILLER_18_1478 VDD VSS sg13g2f_FILL8
XFILLER_18_1486 VDD VSS sg13g2f_FILL8
XFILLER_18_1494 VDD VSS sg13g2f_FILL4
XFILLER_18_1505 VDD VSS sg13g2f_FILL8
XFILLER_18_1513 VDD VSS sg13g2f_FILL8
XFILLER_18_1521 VDD VSS sg13g2f_FILL8
XFILLER_18_1529 VDD VSS sg13g2f_FILL8
XFILLER_18_1537 VDD VSS sg13g2f_FILL8
XFILLER_18_1545 VDD VSS sg13g2f_FILL4
XFILLER_18_1549 VDD VSS sg13g2f_FILL2
XFILLER_19_1390 VDD VSS sg13g2f_FILL8
XFILLER_19_1398 VDD VSS sg13g2f_FILL8
XFILLER_19_1406 VDD VSS sg13g2f_FILL8
XFILLER_19_1414 VDD VSS sg13g2f_FILL8
XFILLER_19_1422 VDD VSS sg13g2f_FILL8
XFILLER_19_1430 VDD VSS sg13g2f_FILL8
XFILLER_19_1438 VDD VSS sg13g2f_FILL8
XFILLER_19_1446 VDD VSS sg13g2f_FILL8
XFILLER_19_1454 VDD VSS sg13g2f_FILL8
XFILLER_19_1462 VDD VSS sg13g2f_FILL8
XFILLER_19_1470 VDD VSS sg13g2f_FILL8
XFILLER_19_1478 VDD VSS sg13g2f_FILL8
XFILLER_19_1486 VDD VSS sg13g2f_FILL8
XFILLER_19_1494 VDD VSS sg13g2f_FILL1
XFILLER_19_1530 VDD VSS sg13g2f_FILL8
XFILLER_19_1538 VDD VSS sg13g2f_FILL8
XFILLER_19_1546 VDD VSS sg13g2f_FILL4
XFILLER_19_1550 VDD VSS sg13g2f_FILL1
XFILLER_20_1390 VDD VSS sg13g2f_FILL8
XFILLER_20_1398 VDD VSS sg13g2f_FILL8
XFILLER_20_1406 VDD VSS sg13g2f_FILL8
XFILLER_20_1414 VDD VSS sg13g2f_FILL8
XFILLER_20_1422 VDD VSS sg13g2f_FILL8
XFILLER_20_1430 VDD VSS sg13g2f_FILL8
XFILLER_20_1438 VDD VSS sg13g2f_FILL8
XFILLER_20_1446 VDD VSS sg13g2f_FILL8
XFILLER_20_1454 VDD VSS sg13g2f_FILL8
XFILLER_20_1462 VDD VSS sg13g2f_FILL8
XFILLER_20_1470 VDD VSS sg13g2f_FILL8
XFILLER_20_1478 VDD VSS sg13g2f_FILL1
XFILLER_20_1505 VDD VSS sg13g2f_FILL2
XFILLER_20_1507 VDD VSS sg13g2f_FILL1
XFILLER_20_1538 VDD VSS sg13g2f_FILL8
XFILLER_20_1546 VDD VSS sg13g2f_FILL4
XFILLER_20_1550 VDD VSS sg13g2f_FILL1
XFILLER_21_1390 VDD VSS sg13g2f_FILL8
XFILLER_21_1398 VDD VSS sg13g2f_FILL8
XFILLER_21_1406 VDD VSS sg13g2f_FILL8
XFILLER_21_1414 VDD VSS sg13g2f_FILL8
XFILLER_21_1422 VDD VSS sg13g2f_FILL8
XFILLER_21_1430 VDD VSS sg13g2f_FILL8
XFILLER_21_1438 VDD VSS sg13g2f_FILL8
XFILLER_21_1446 VDD VSS sg13g2f_FILL8
XFILLER_21_1454 VDD VSS sg13g2f_FILL8
XFILLER_21_1462 VDD VSS sg13g2f_FILL8
XFILLER_21_1470 VDD VSS sg13g2f_FILL8
XFILLER_21_1478 VDD VSS sg13g2f_FILL8
XFILLER_21_1486 VDD VSS sg13g2f_FILL8
XFILLER_21_1494 VDD VSS sg13g2f_FILL8
XFILLER_21_1502 VDD VSS sg13g2f_FILL8
XFILLER_21_1510 VDD VSS sg13g2f_FILL8
XFILLER_21_1518 VDD VSS sg13g2f_FILL8
XFILLER_21_1526 VDD VSS sg13g2f_FILL8
XFILLER_21_1534 VDD VSS sg13g2f_FILL8
XFILLER_21_1542 VDD VSS sg13g2f_FILL8
XFILLER_21_1550 VDD VSS sg13g2f_FILL1
XFILLER_22_7 AVDD VSS sg13g2f_FILL4
XFILLER_22_11 AVDD VSS sg13g2f_FILL1
XFILLER_22_47 AVDD VSS sg13g2f_FILL1
XFILLER_22_119 AVDD VSS sg13g2f_FILL8
XFILLER_22_127 AVDD VSS sg13g2f_FILL8
XFILLER_22_135 AVDD VSS sg13g2f_FILL8
XFILLER_22_143 AVDD VSS sg13g2f_FILL8
XFILLER_22_151 AVDD VSS sg13g2f_FILL8
XFILLER_22_159 AVDD VSS sg13g2f_FILL8
XFILLER_22_167 AVDD VSS sg13g2f_FILL8
XFILLER_22_175 AVDD VSS sg13g2f_FILL8
XFILLER_22_183 AVDD VSS sg13g2f_FILL8
XFILLER_22_191 AVDD VSS sg13g2f_FILL8
XFILLER_22_199 AVDD VSS sg13g2f_FILL8
XFILLER_22_207 AVDD VSS sg13g2f_FILL8
XFILLER_22_215 AVDD VSS sg13g2f_FILL8
XFILLER_22_223 AVDD VSS sg13g2f_FILL1
XFILLER_22_231 AVDD VSS sg13g2f_FILL8
XFILLER_22_239 AVDD VSS sg13g2f_FILL8
XFILLER_22_247 AVDD VSS sg13g2f_FILL8
XFILLER_22_255 AVDD VSS sg13g2f_FILL8
XFILLER_22_263 AVDD VSS sg13g2f_FILL8
XFILLER_22_271 AVDD VSS sg13g2f_FILL8
XFILLER_22_279 AVDD VSS sg13g2f_FILL8
XFILLER_22_287 AVDD VSS sg13g2f_FILL8
XFILLER_22_295 AVDD VSS sg13g2f_FILL8
XFILLER_22_303 AVDD VSS sg13g2f_FILL8
XFILLER_22_311 AVDD VSS sg13g2f_FILL8
XFILLER_22_319 AVDD VSS sg13g2f_FILL8
XFILLER_22_327 AVDD VSS sg13g2f_FILL8
XFILLER_22_335 AVDD VSS sg13g2f_FILL1
XFILLER_22_343 AVDD VSS sg13g2f_FILL8
XFILLER_22_351 AVDD VSS sg13g2f_FILL8
XFILLER_22_359 AVDD VSS sg13g2f_FILL8
XFILLER_22_367 AVDD VSS sg13g2f_FILL8
XFILLER_22_375 AVDD VSS sg13g2f_FILL8
XFILLER_22_383 AVDD VSS sg13g2f_FILL1
XFILLER_22_455 AVDD VSS sg13g2f_FILL8
XFILLER_22_463 AVDD VSS sg13g2f_FILL8
XFILLER_22_471 AVDD VSS sg13g2f_FILL8
XFILLER_22_479 AVDD VSS sg13g2f_FILL8
XFILLER_22_487 AVDD VSS sg13g2f_FILL8
XFILLER_22_495 AVDD VSS sg13g2f_FILL8
XFILLER_22_503 AVDD VSS sg13g2f_FILL8
XFILLER_22_511 AVDD VSS sg13g2f_FILL8
XFILLER_22_519 AVDD VSS sg13g2f_FILL8
XFILLER_22_527 AVDD VSS sg13g2f_FILL8
XFILLER_22_535 AVDD VSS sg13g2f_FILL8
XFILLER_22_543 AVDD VSS sg13g2f_FILL8
XFILLER_22_551 AVDD VSS sg13g2f_FILL8
XFILLER_22_559 AVDD VSS sg13g2f_FILL1
XFILLER_22_567 AVDD VSS sg13g2f_FILL8
XFILLER_22_575 AVDD VSS sg13g2f_FILL8
XFILLER_22_583 AVDD VSS sg13g2f_FILL8
XFILLER_22_591 AVDD VSS sg13g2f_FILL8
XFILLER_22_599 AVDD VSS sg13g2f_FILL8
XFILLER_22_607 AVDD VSS sg13g2f_FILL8
XFILLER_22_615 AVDD VSS sg13g2f_FILL8
XFILLER_22_623 AVDD VSS sg13g2f_FILL8
XFILLER_22_631 AVDD VSS sg13g2f_FILL8
XFILLER_22_639 AVDD VSS sg13g2f_FILL8
XFILLER_22_647 AVDD VSS sg13g2f_FILL8
XFILLER_22_655 AVDD VSS sg13g2f_FILL8
XFILLER_22_663 AVDD VSS sg13g2f_FILL8
XFILLER_22_671 AVDD VSS sg13g2f_FILL1
XFILLER_22_679 AVDD VSS sg13g2f_FILL8
XFILLER_22_687 AVDD VSS sg13g2f_FILL8
XFILLER_22_695 AVDD VSS sg13g2f_FILL8
XFILLER_22_703 AVDD VSS sg13g2f_FILL8
XFILLER_22_711 AVDD VSS sg13g2f_FILL8
XFILLER_22_719 AVDD VSS sg13g2f_FILL8
XFILLER_22_727 AVDD VSS sg13g2f_FILL8
XFILLER_22_735 AVDD VSS sg13g2f_FILL8
XFILLER_22_743 AVDD VSS sg13g2f_FILL8
XFILLER_22_751 AVDD VSS sg13g2f_FILL8
XFILLER_22_759 AVDD VSS sg13g2f_FILL8
XFILLER_22_767 AVDD VSS sg13g2f_FILL8
XFILLER_22_775 AVDD VSS sg13g2f_FILL8
XFILLER_22_783 AVDD VSS sg13g2f_FILL1
XFILLER_22_791 AVDD VSS sg13g2f_FILL8
XFILLER_22_799 AVDD VSS sg13g2f_FILL8
XFILLER_22_807 AVDD VSS sg13g2f_FILL8
XFILLER_22_815 AVDD VSS sg13g2f_FILL8
XFILLER_22_823 AVDD VSS sg13g2f_FILL8
XFILLER_22_831 AVDD VSS sg13g2f_FILL8
XFILLER_22_839 AVDD VSS sg13g2f_FILL8
XFILLER_22_847 AVDD VSS sg13g2f_FILL8
XFILLER_22_855 AVDD VSS sg13g2f_FILL8
XFILLER_22_863 AVDD VSS sg13g2f_FILL8
XFILLER_22_871 AVDD VSS sg13g2f_FILL8
XFILLER_22_879 AVDD VSS sg13g2f_FILL8
XFILLER_22_887 AVDD VSS sg13g2f_FILL8
XFILLER_22_895 AVDD VSS sg13g2f_FILL1
XFILLER_22_903 AVDD VSS sg13g2f_FILL8
XFILLER_22_911 AVDD VSS sg13g2f_FILL8
XFILLER_22_919 AVDD VSS sg13g2f_FILL8
XFILLER_22_927 AVDD VSS sg13g2f_FILL8
XFILLER_22_935 AVDD VSS sg13g2f_FILL8
XFILLER_22_943 AVDD VSS sg13g2f_FILL8
XFILLER_22_951 AVDD VSS sg13g2f_FILL8
XFILLER_22_959 AVDD VSS sg13g2f_FILL8
XFILLER_22_967 AVDD VSS sg13g2f_FILL8
XFILLER_22_975 AVDD VSS sg13g2f_FILL8
XFILLER_22_983 AVDD VSS sg13g2f_FILL8
XFILLER_22_991 AVDD VSS sg13g2f_FILL8
XFILLER_22_999 AVDD VSS sg13g2f_FILL8
XFILLER_22_1007 AVDD VSS sg13g2f_FILL1
XFILLER_22_1015 AVDD VSS sg13g2f_FILL8
XFILLER_22_1023 AVDD VSS sg13g2f_FILL8
XFILLER_22_1031 AVDD VSS sg13g2f_FILL8
XFILLER_22_1039 AVDD VSS sg13g2f_FILL8
XFILLER_22_1047 AVDD VSS sg13g2f_FILL8
XFILLER_22_1055 AVDD VSS sg13g2f_FILL8
XFILLER_22_1063 AVDD VSS sg13g2f_FILL8
XFILLER_22_1071 AVDD VSS sg13g2f_FILL8
XFILLER_22_1079 AVDD VSS sg13g2f_FILL8
XFILLER_22_1087 AVDD VSS sg13g2f_FILL8
XFILLER_22_1095 AVDD VSS sg13g2f_FILL8
XFILLER_22_1103 AVDD VSS sg13g2f_FILL8
XFILLER_22_1111 AVDD VSS sg13g2f_FILL8
XFILLER_22_1119 AVDD VSS sg13g2f_FILL1
XFILLER_22_1127 AVDD VSS sg13g2f_FILL8
XFILLER_22_1135 AVDD VSS sg13g2f_FILL4
XFILLER_22_1139 AVDD VSS sg13g2f_FILL2
XFILLER_22_1152 AVDD VSS sg13g2f_FILL8
XFILLER_22_1160 AVDD VSS sg13g2f_FILL8
XFILLER_22_1168 AVDD VSS sg13g2f_FILL8
XFILLER_22_1176 AVDD VSS sg13g2f_FILL8
XFILLER_22_1184 AVDD VSS sg13g2f_FILL8
XFILLER_22_1192 AVDD VSS sg13g2f_FILL8
XFILLER_22_1200 AVDD VSS sg13g2f_FILL8
XFILLER_22_1208 AVDD VSS sg13g2f_FILL8
XFILLER_22_1216 AVDD VSS sg13g2f_FILL8
XFILLER_22_1224 AVDD VSS sg13g2f_FILL8
XFILLER_22_1239 AVDD VSS sg13g2f_FILL8
XFILLER_22_1247 AVDD VSS sg13g2f_FILL8
XFILLER_22_1255 AVDD VSS sg13g2f_FILL8
XFILLER_22_1263 AVDD VSS sg13g2f_FILL4
XFILLER_22_1267 AVDD VSS sg13g2f_FILL1
XFILLER_22_1390 VDD VSS sg13g2f_FILL8
XFILLER_22_1398 VDD VSS sg13g2f_FILL8
XFILLER_22_1406 VDD VSS sg13g2f_FILL8
XFILLER_22_1414 VDD VSS sg13g2f_FILL8
XFILLER_22_1422 VDD VSS sg13g2f_FILL8
XFILLER_22_1430 VDD VSS sg13g2f_FILL8
XFILLER_22_1438 VDD VSS sg13g2f_FILL8
XFILLER_22_1446 VDD VSS sg13g2f_FILL8
XFILLER_22_1454 VDD VSS sg13g2f_FILL8
XFILLER_22_1462 VDD VSS sg13g2f_FILL8
XFILLER_22_1470 VDD VSS sg13g2f_FILL8
XFILLER_22_1478 VDD VSS sg13g2f_FILL8
XFILLER_22_1486 VDD VSS sg13g2f_FILL8
XFILLER_22_1494 VDD VSS sg13g2f_FILL4
XFILLER_22_1547 VDD VSS sg13g2f_FILL4
XFILLER_23_7 AVDD VSS sg13g2f_FILL4
XFILLER_23_11 AVDD VSS sg13g2f_FILL1
XFILLER_23_58 AVDD VSS sg13g2f_FILL4
XFILLER_23_126 AVDD VSS sg13g2f_FILL8
XFILLER_23_134 AVDD VSS sg13g2f_FILL8
XFILLER_23_142 AVDD VSS sg13g2f_FILL8
XFILLER_23_150 AVDD VSS sg13g2f_FILL8
XFILLER_23_158 AVDD VSS sg13g2f_FILL8
XFILLER_23_166 AVDD VSS sg13g2f_FILL8
XFILLER_23_174 AVDD VSS sg13g2f_FILL8
XFILLER_23_182 AVDD VSS sg13g2f_FILL8
XFILLER_23_190 AVDD VSS sg13g2f_FILL8
XFILLER_23_198 AVDD VSS sg13g2f_FILL8
XFILLER_23_206 AVDD VSS sg13g2f_FILL8
XFILLER_23_214 AVDD VSS sg13g2f_FILL8
XFILLER_23_222 AVDD VSS sg13g2f_FILL8
XFILLER_23_230 AVDD VSS sg13g2f_FILL1
XFILLER_23_238 AVDD VSS sg13g2f_FILL8
XFILLER_23_246 AVDD VSS sg13g2f_FILL8
XFILLER_23_254 AVDD VSS sg13g2f_FILL8
XFILLER_23_262 AVDD VSS sg13g2f_FILL8
XFILLER_23_270 AVDD VSS sg13g2f_FILL8
XFILLER_23_278 AVDD VSS sg13g2f_FILL8
XFILLER_23_286 AVDD VSS sg13g2f_FILL8
XFILLER_23_294 AVDD VSS sg13g2f_FILL8
XFILLER_23_302 AVDD VSS sg13g2f_FILL8
XFILLER_23_310 AVDD VSS sg13g2f_FILL8
XFILLER_23_318 AVDD VSS sg13g2f_FILL8
XFILLER_23_326 AVDD VSS sg13g2f_FILL8
XFILLER_23_334 AVDD VSS sg13g2f_FILL8
XFILLER_23_342 AVDD VSS sg13g2f_FILL8
XFILLER_23_350 AVDD VSS sg13g2f_FILL8
XFILLER_23_358 AVDD VSS sg13g2f_FILL8
XFILLER_23_366 AVDD VSS sg13g2f_FILL8
XFILLER_23_374 AVDD VSS sg13g2f_FILL8
XFILLER_23_382 AVDD VSS sg13g2f_FILL8
XFILLER_23_390 AVDD VSS sg13g2f_FILL4
XFILLER_23_394 AVDD VSS sg13g2f_FILL1
XFILLER_23_459 AVDD VSS sg13g2f_FILL2
XFILLER_23_461 AVDD VSS sg13g2f_FILL1
XFILLER_23_469 AVDD VSS sg13g2f_FILL8
XFILLER_23_477 AVDD VSS sg13g2f_FILL8
XFILLER_23_485 AVDD VSS sg13g2f_FILL8
XFILLER_23_493 AVDD VSS sg13g2f_FILL8
XFILLER_23_501 AVDD VSS sg13g2f_FILL8
XFILLER_23_509 AVDD VSS sg13g2f_FILL8
XFILLER_23_517 AVDD VSS sg13g2f_FILL8
XFILLER_23_525 AVDD VSS sg13g2f_FILL8
XFILLER_23_533 AVDD VSS sg13g2f_FILL8
XFILLER_23_541 AVDD VSS sg13g2f_FILL8
XFILLER_23_549 AVDD VSS sg13g2f_FILL8
XFILLER_23_557 AVDD VSS sg13g2f_FILL1
XFILLER_23_622 AVDD VSS sg13g2f_FILL8
XFILLER_23_630 AVDD VSS sg13g2f_FILL8
XFILLER_23_638 AVDD VSS sg13g2f_FILL8
XFILLER_23_646 AVDD VSS sg13g2f_FILL8
XFILLER_23_654 AVDD VSS sg13g2f_FILL8
XFILLER_23_662 AVDD VSS sg13g2f_FILL8
XFILLER_23_670 AVDD VSS sg13g2f_FILL8
XFILLER_23_678 AVDD VSS sg13g2f_FILL8
XFILLER_23_686 AVDD VSS sg13g2f_FILL4
XFILLER_23_690 AVDD VSS sg13g2f_FILL2
XFILLER_23_692 AVDD VSS sg13g2f_FILL1
XFILLER_23_700 AVDD VSS sg13g2f_FILL8
XFILLER_23_708 AVDD VSS sg13g2f_FILL8
XFILLER_23_716 AVDD VSS sg13g2f_FILL8
XFILLER_23_724 AVDD VSS sg13g2f_FILL8
XFILLER_23_732 AVDD VSS sg13g2f_FILL8
XFILLER_23_740 AVDD VSS sg13g2f_FILL8
XFILLER_23_748 AVDD VSS sg13g2f_FILL8
XFILLER_23_756 AVDD VSS sg13g2f_FILL8
XFILLER_23_764 AVDD VSS sg13g2f_FILL8
XFILLER_23_772 AVDD VSS sg13g2f_FILL8
XFILLER_23_780 AVDD VSS sg13g2f_FILL8
XFILLER_23_788 AVDD VSS sg13g2f_FILL8
XFILLER_23_796 AVDD VSS sg13g2f_FILL8
XFILLER_23_804 AVDD VSS sg13g2f_FILL8
XFILLER_23_812 AVDD VSS sg13g2f_FILL8
XFILLER_23_820 AVDD VSS sg13g2f_FILL8
XFILLER_23_828 AVDD VSS sg13g2f_FILL8
XFILLER_23_836 AVDD VSS sg13g2f_FILL8
XFILLER_23_844 AVDD VSS sg13g2f_FILL8
XFILLER_23_868 AVDD VSS sg13g2f_FILL8
XFILLER_23_876 AVDD VSS sg13g2f_FILL4
XFILLER_23_905 AVDD VSS sg13g2f_FILL8
XFILLER_23_913 AVDD VSS sg13g2f_FILL8
XFILLER_23_921 AVDD VSS sg13g2f_FILL2
XFILLER_23_923 AVDD VSS sg13g2f_FILL1
XFILLER_23_931 AVDD VSS sg13g2f_FILL8
XFILLER_23_939 AVDD VSS sg13g2f_FILL8
XFILLER_23_947 AVDD VSS sg13g2f_FILL8
XFILLER_23_955 AVDD VSS sg13g2f_FILL8
XFILLER_23_963 AVDD VSS sg13g2f_FILL8
XFILLER_23_971 AVDD VSS sg13g2f_FILL8
XFILLER_23_979 AVDD VSS sg13g2f_FILL8
XFILLER_23_987 AVDD VSS sg13g2f_FILL8
XFILLER_23_995 AVDD VSS sg13g2f_FILL8
XFILLER_23_1003 AVDD VSS sg13g2f_FILL8
XFILLER_23_1011 AVDD VSS sg13g2f_FILL8
XFILLER_23_1019 AVDD VSS sg13g2f_FILL2
XFILLER_23_1021 AVDD VSS sg13g2f_FILL1
XFILLER_23_1038 AVDD VSS sg13g2f_FILL8
XFILLER_23_1110 AVDD VSS sg13g2f_FILL8
XFILLER_23_1118 AVDD VSS sg13g2f_FILL8
XFILLER_23_1126 AVDD VSS sg13g2f_FILL8
XFILLER_23_1150 AVDD VSS sg13g2f_FILL4
XFILLER_23_1154 AVDD VSS sg13g2f_FILL1
XFILLER_23_1162 AVDD VSS sg13g2f_FILL8
XFILLER_23_1170 AVDD VSS sg13g2f_FILL8
XFILLER_23_1178 AVDD VSS sg13g2f_FILL8
XFILLER_23_1186 AVDD VSS sg13g2f_FILL8
XFILLER_23_1194 AVDD VSS sg13g2f_FILL8
XFILLER_23_1202 AVDD VSS sg13g2f_FILL8
XFILLER_23_1210 AVDD VSS sg13g2f_FILL8
XFILLER_23_1218 AVDD VSS sg13g2f_FILL8
XFILLER_23_1226 AVDD VSS sg13g2f_FILL8
XFILLER_23_1234 AVDD VSS sg13g2f_FILL8
XFILLER_23_1242 AVDD VSS sg13g2f_FILL8
XFILLER_23_1250 AVDD VSS sg13g2f_FILL8
XFILLER_23_1258 AVDD VSS sg13g2f_FILL8
XFILLER_23_1266 AVDD VSS sg13g2f_FILL2
XFILLER_23_1390 VDD VSS sg13g2f_FILL8
XFILLER_23_1398 VDD VSS sg13g2f_FILL8
XFILLER_23_1406 VDD VSS sg13g2f_FILL8
XFILLER_23_1414 VDD VSS sg13g2f_FILL8
XFILLER_23_1422 VDD VSS sg13g2f_FILL8
XFILLER_23_1430 VDD VSS sg13g2f_FILL8
XFILLER_23_1438 VDD VSS sg13g2f_FILL8
XFILLER_23_1446 VDD VSS sg13g2f_FILL8
XFILLER_23_1454 VDD VSS sg13g2f_FILL8
XFILLER_23_1462 VDD VSS sg13g2f_FILL8
XFILLER_23_1470 VDD VSS sg13g2f_FILL8
XFILLER_23_1478 VDD VSS sg13g2f_FILL8
XFILLER_23_1486 VDD VSS sg13g2f_FILL8
XFILLER_23_1494 VDD VSS sg13g2f_FILL8
XFILLER_23_1502 VDD VSS sg13g2f_FILL1
XFILLER_23_1545 VDD VSS sg13g2f_FILL4
XFILLER_23_1549 VDD VSS sg13g2f_FILL2
XFILLER_24_7 AVDD VSS sg13g2f_FILL4
XFILLER_24_11 AVDD VSS sg13g2f_FILL1
XFILLER_24_119 AVDD VSS sg13g2f_FILL8
XFILLER_24_127 AVDD VSS sg13g2f_FILL8
XFILLER_24_135 AVDD VSS sg13g2f_FILL8
XFILLER_24_143 AVDD VSS sg13g2f_FILL8
XFILLER_24_151 AVDD VSS sg13g2f_FILL8
XFILLER_24_159 AVDD VSS sg13g2f_FILL8
XFILLER_24_167 AVDD VSS sg13g2f_FILL8
XFILLER_24_175 AVDD VSS sg13g2f_FILL8
XFILLER_24_183 AVDD VSS sg13g2f_FILL8
XFILLER_24_191 AVDD VSS sg13g2f_FILL8
XFILLER_24_199 AVDD VSS sg13g2f_FILL8
XFILLER_24_207 AVDD VSS sg13g2f_FILL8
XFILLER_24_215 AVDD VSS sg13g2f_FILL8
XFILLER_24_223 AVDD VSS sg13g2f_FILL1
XFILLER_24_247 AVDD VSS sg13g2f_FILL8
XFILLER_24_255 AVDD VSS sg13g2f_FILL8
XFILLER_24_263 AVDD VSS sg13g2f_FILL8
XFILLER_24_271 AVDD VSS sg13g2f_FILL8
XFILLER_24_279 AVDD VSS sg13g2f_FILL8
XFILLER_24_287 AVDD VSS sg13g2f_FILL8
XFILLER_24_295 AVDD VSS sg13g2f_FILL8
XFILLER_24_303 AVDD VSS sg13g2f_FILL8
XFILLER_24_311 AVDD VSS sg13g2f_FILL8
XFILLER_24_319 AVDD VSS sg13g2f_FILL8
XFILLER_24_327 AVDD VSS sg13g2f_FILL8
XFILLER_24_335 AVDD VSS sg13g2f_FILL1
XFILLER_24_343 AVDD VSS sg13g2f_FILL8
XFILLER_24_351 AVDD VSS sg13g2f_FILL1
XFILLER_24_374 AVDD VSS sg13g2f_FILL8
XFILLER_24_382 AVDD VSS sg13g2f_FILL2
XFILLER_24_455 AVDD VSS sg13g2f_FILL8
XFILLER_24_463 AVDD VSS sg13g2f_FILL8
XFILLER_24_471 AVDD VSS sg13g2f_FILL8
XFILLER_24_479 AVDD VSS sg13g2f_FILL8
XFILLER_24_487 AVDD VSS sg13g2f_FILL8
XFILLER_24_495 AVDD VSS sg13g2f_FILL8
XFILLER_24_503 AVDD VSS sg13g2f_FILL8
XFILLER_24_511 AVDD VSS sg13g2f_FILL8
XFILLER_24_519 AVDD VSS sg13g2f_FILL8
XFILLER_24_527 AVDD VSS sg13g2f_FILL8
XFILLER_24_535 AVDD VSS sg13g2f_FILL8
XFILLER_24_543 AVDD VSS sg13g2f_FILL8
XFILLER_24_551 AVDD VSS sg13g2f_FILL8
XFILLER_24_559 AVDD VSS sg13g2f_FILL1
XFILLER_24_567 AVDD VSS sg13g2f_FILL8
XFILLER_24_575 AVDD VSS sg13g2f_FILL8
XFILLER_24_583 AVDD VSS sg13g2f_FILL8
XFILLER_24_591 AVDD VSS sg13g2f_FILL8
XFILLER_24_599 AVDD VSS sg13g2f_FILL8
XFILLER_24_607 AVDD VSS sg13g2f_FILL8
XFILLER_24_615 AVDD VSS sg13g2f_FILL8
XFILLER_24_623 AVDD VSS sg13g2f_FILL8
XFILLER_24_631 AVDD VSS sg13g2f_FILL8
XFILLER_24_639 AVDD VSS sg13g2f_FILL8
XFILLER_24_647 AVDD VSS sg13g2f_FILL8
XFILLER_24_655 AVDD VSS sg13g2f_FILL8
XFILLER_24_663 AVDD VSS sg13g2f_FILL8
XFILLER_24_671 AVDD VSS sg13g2f_FILL1
XFILLER_24_679 AVDD VSS sg13g2f_FILL2
XFILLER_24_681 AVDD VSS sg13g2f_FILL1
XFILLER_24_746 AVDD VSS sg13g2f_FILL8
XFILLER_24_754 AVDD VSS sg13g2f_FILL8
XFILLER_24_762 AVDD VSS sg13g2f_FILL8
XFILLER_24_770 AVDD VSS sg13g2f_FILL8
XFILLER_24_778 AVDD VSS sg13g2f_FILL4
XFILLER_24_782 AVDD VSS sg13g2f_FILL2
XFILLER_24_855 AVDD VSS sg13g2f_FILL8
XFILLER_24_863 AVDD VSS sg13g2f_FILL8
XFILLER_24_871 AVDD VSS sg13g2f_FILL8
XFILLER_24_879 AVDD VSS sg13g2f_FILL1
XFILLER_24_928 AVDD VSS sg13g2f_FILL2
XFILLER_24_994 AVDD VSS sg13g2f_FILL8
XFILLER_24_1002 AVDD VSS sg13g2f_FILL4
XFILLER_24_1006 AVDD VSS sg13g2f_FILL2
XFILLER_24_1101 AVDD VSS sg13g2f_FILL4
XFILLER_24_1105 AVDD VSS sg13g2f_FILL2
XFILLER_24_1118 AVDD VSS sg13g2f_FILL2
XFILLER_24_1127 AVDD VSS sg13g2f_FILL1
XFILLER_24_1153 AVDD VSS sg13g2f_FILL4
XFILLER_24_1198 AVDD VSS sg13g2f_FILL8
XFILLER_24_1206 AVDD VSS sg13g2f_FILL8
XFILLER_24_1214 AVDD VSS sg13g2f_FILL8
XFILLER_24_1222 AVDD VSS sg13g2f_FILL8
XFILLER_24_1230 AVDD VSS sg13g2f_FILL2
XFILLER_24_1239 AVDD VSS sg13g2f_FILL8
XFILLER_24_1247 AVDD VSS sg13g2f_FILL8
XFILLER_24_1255 AVDD VSS sg13g2f_FILL8
XFILLER_24_1263 AVDD VSS sg13g2f_FILL4
XFILLER_24_1267 AVDD VSS sg13g2f_FILL1
XFILLER_24_1398 VDD VSS sg13g2f_FILL8
XFILLER_24_1406 VDD VSS sg13g2f_FILL8
XFILLER_24_1414 VDD VSS sg13g2f_FILL8
XFILLER_24_1422 VDD VSS sg13g2f_FILL8
XFILLER_24_1430 VDD VSS sg13g2f_FILL8
XFILLER_24_1438 VDD VSS sg13g2f_FILL8
XFILLER_24_1446 VDD VSS sg13g2f_FILL8
XFILLER_24_1454 VDD VSS sg13g2f_FILL8
XFILLER_24_1462 VDD VSS sg13g2f_FILL8
XFILLER_24_1470 VDD VSS sg13g2f_FILL8
XFILLER_24_1478 VDD VSS sg13g2f_FILL8
XFILLER_24_1486 VDD VSS sg13g2f_FILL8
XFILLER_24_1494 VDD VSS sg13g2f_FILL4
XFILLER_24_1513 VDD VSS sg13g2f_FILL8
XFILLER_24_1521 VDD VSS sg13g2f_FILL8
XFILLER_24_1529 VDD VSS sg13g2f_FILL8
XFILLER_24_1537 VDD VSS sg13g2f_FILL8
XFILLER_24_1545 VDD VSS sg13g2f_FILL4
XFILLER_24_1549 VDD VSS sg13g2f_FILL2
XFILLER_25_151 AVDD VSS sg13g2f_FILL8
XFILLER_25_159 AVDD VSS sg13g2f_FILL8
XFILLER_25_167 AVDD VSS sg13g2f_FILL8
XFILLER_25_175 AVDD VSS sg13g2f_FILL4
XFILLER_25_179 AVDD VSS sg13g2f_FILL1
XFILLER_25_205 AVDD VSS sg13g2f_FILL8
XFILLER_25_238 AVDD VSS sg13g2f_FILL8
XFILLER_25_246 AVDD VSS sg13g2f_FILL8
XFILLER_25_254 AVDD VSS sg13g2f_FILL8
XFILLER_25_262 AVDD VSS sg13g2f_FILL2
XFILLER_25_289 AVDD VSS sg13g2f_FILL8
XFILLER_25_297 AVDD VSS sg13g2f_FILL8
XFILLER_25_305 AVDD VSS sg13g2f_FILL8
XFILLER_25_313 AVDD VSS sg13g2f_FILL4
XFILLER_25_317 AVDD VSS sg13g2f_FILL2
XFILLER_25_319 AVDD VSS sg13g2f_FILL1
XFILLER_25_336 AVDD VSS sg13g2f_FILL2
XFILLER_25_368 AVDD VSS sg13g2f_FILL4
XFILLER_25_372 AVDD VSS sg13g2f_FILL2
XFILLER_25_374 AVDD VSS sg13g2f_FILL1
XFILLER_25_382 AVDD VSS sg13g2f_FILL2
XFILLER_25_427 AVDD VSS sg13g2f_FILL4
XFILLER_25_431 AVDD VSS sg13g2f_FILL2
XFILLER_25_433 AVDD VSS sg13g2f_FILL1
XFILLER_25_498 AVDD VSS sg13g2f_FILL8
XFILLER_25_506 AVDD VSS sg13g2f_FILL8
XFILLER_25_514 AVDD VSS sg13g2f_FILL8
XFILLER_25_522 AVDD VSS sg13g2f_FILL8
XFILLER_25_530 AVDD VSS sg13g2f_FILL8
XFILLER_25_538 AVDD VSS sg13g2f_FILL2
XFILLER_25_540 AVDD VSS sg13g2f_FILL1
XFILLER_25_605 AVDD VSS sg13g2f_FILL1
XFILLER_25_613 AVDD VSS sg13g2f_FILL8
XFILLER_25_621 AVDD VSS sg13g2f_FILL8
XFILLER_25_629 AVDD VSS sg13g2f_FILL2
XFILLER_25_631 AVDD VSS sg13g2f_FILL1
XFILLER_25_665 AVDD VSS sg13g2f_FILL8
XFILLER_25_673 AVDD VSS sg13g2f_FILL2
XFILLER_25_675 AVDD VSS sg13g2f_FILL1
XFILLER_25_740 AVDD VSS sg13g2f_FILL8
XFILLER_25_748 AVDD VSS sg13g2f_FILL8
XFILLER_25_820 AVDD VSS sg13g2f_FILL1
XFILLER_25_844 AVDD VSS sg13g2f_FILL1
XFILLER_25_870 AVDD VSS sg13g2f_FILL8
XFILLER_25_878 AVDD VSS sg13g2f_FILL2
XFILLER_25_960 AVDD VSS sg13g2f_FILL4
XFILLER_25_964 AVDD VSS sg13g2f_FILL1
XFILLER_25_986 AVDD VSS sg13g2f_FILL8
XFILLER_25_994 AVDD VSS sg13g2f_FILL8
XFILLER_25_1002 AVDD VSS sg13g2f_FILL8
XFILLER_25_1010 AVDD VSS sg13g2f_FILL4
XFILLER_25_1014 AVDD VSS sg13g2f_FILL2
XFILLER_25_1041 AVDD VSS sg13g2f_FILL2
XFILLER_25_1116 AVDD VSS sg13g2f_FILL8
XFILLER_25_1124 AVDD VSS sg13g2f_FILL4
XFILLER_25_1139 AVDD VSS sg13g2f_FILL2
XFILLER_25_1141 AVDD VSS sg13g2f_FILL1
XFILLER_25_1206 AVDD VSS sg13g2f_FILL8
XFILLER_25_1214 AVDD VSS sg13g2f_FILL8
XFILLER_25_1222 AVDD VSS sg13g2f_FILL8
XFILLER_25_1230 AVDD VSS sg13g2f_FILL8
XFILLER_25_1238 AVDD VSS sg13g2f_FILL8
XFILLER_25_1246 AVDD VSS sg13g2f_FILL8
XFILLER_25_1254 AVDD VSS sg13g2f_FILL8
XFILLER_25_1262 AVDD VSS sg13g2f_FILL4
XFILLER_25_1266 AVDD VSS sg13g2f_FILL2
XFILLER_25_1390 VDD VSS sg13g2f_FILL8
XFILLER_25_1398 VDD VSS sg13g2f_FILL8
XFILLER_25_1406 VDD VSS sg13g2f_FILL8
XFILLER_25_1414 VDD VSS sg13g2f_FILL8
XFILLER_25_1422 VDD VSS sg13g2f_FILL8
XFILLER_25_1430 VDD VSS sg13g2f_FILL8
XFILLER_25_1438 VDD VSS sg13g2f_FILL8
XFILLER_25_1446 VDD VSS sg13g2f_FILL8
XFILLER_25_1454 VDD VSS sg13g2f_FILL8
XFILLER_25_1462 VDD VSS sg13g2f_FILL8
XFILLER_25_1470 VDD VSS sg13g2f_FILL8
XFILLER_25_1478 VDD VSS sg13g2f_FILL8
XFILLER_25_1486 VDD VSS sg13g2f_FILL8
XFILLER_25_1494 VDD VSS sg13g2f_FILL8
XFILLER_25_1502 VDD VSS sg13g2f_FILL8
XFILLER_25_1510 VDD VSS sg13g2f_FILL4
XFILLER_25_1514 VDD VSS sg13g2f_FILL2
XFILLER_25_1535 VDD VSS sg13g2f_FILL8
XFILLER_25_1543 VDD VSS sg13g2f_FILL8
XFILLER_26_405 AVDD VSS sg13g2f_FILL4
XFILLER_26_409 AVDD VSS sg13g2f_FILL1
XFILLER_26_497 AVDD VSS sg13g2f_FILL8
XFILLER_26_505 AVDD VSS sg13g2f_FILL2
XFILLER_26_507 AVDD VSS sg13g2f_FILL1
XFILLER_26_524 AVDD VSS sg13g2f_FILL8
XFILLER_26_532 AVDD VSS sg13g2f_FILL1
XFILLER_26_622 AVDD VSS sg13g2f_FILL8
XFILLER_26_630 AVDD VSS sg13g2f_FILL8
XFILLER_26_638 AVDD VSS sg13g2f_FILL2
XFILLER_26_656 AVDD VSS sg13g2f_FILL1
XFILLER_26_744 AVDD VSS sg13g2f_FILL8
XFILLER_26_752 AVDD VSS sg13g2f_FILL4
XFILLER_26_772 AVDD VSS sg13g2f_FILL1
XFILLER_26_846 AVDD VSS sg13g2f_FILL4
XFILLER_26_850 AVDD VSS sg13g2f_FILL1
XFILLER_26_870 AVDD VSS sg13g2f_FILL8
XFILLER_26_878 AVDD VSS sg13g2f_FILL2
XFILLER_26_937 AVDD VSS sg13g2f_FILL4
XFILLER_26_970 AVDD VSS sg13g2f_FILL8
XFILLER_26_994 AVDD VSS sg13g2f_FILL8
XFILLER_26_1002 AVDD VSS sg13g2f_FILL8
XFILLER_26_1010 AVDD VSS sg13g2f_FILL8
XFILLER_26_1099 AVDD VSS sg13g2f_FILL8
XFILLER_26_1107 AVDD VSS sg13g2f_FILL8
XFILLER_26_1115 AVDD VSS sg13g2f_FILL8
XFILLER_26_1123 AVDD VSS sg13g2f_FILL8
XFILLER_26_1131 AVDD VSS sg13g2f_FILL4
XFILLER_26_1135 AVDD VSS sg13g2f_FILL2
XFILLER_26_1162 AVDD VSS sg13g2f_FILL2
XFILLER_26_1190 AVDD VSS sg13g2f_FILL8
XFILLER_26_1198 AVDD VSS sg13g2f_FILL4
XFILLER_26_1202 AVDD VSS sg13g2f_FILL2
XFILLER_26_1406 VDD VSS sg13g2f_FILL8
XFILLER_26_1414 VDD VSS sg13g2f_FILL8
XFILLER_26_1422 VDD VSS sg13g2f_FILL8
XFILLER_26_1430 VDD VSS sg13g2f_FILL8
XFILLER_26_1438 VDD VSS sg13g2f_FILL8
XFILLER_26_1446 VDD VSS sg13g2f_FILL8
XFILLER_26_1454 VDD VSS sg13g2f_FILL8
XFILLER_26_1462 VDD VSS sg13g2f_FILL8
XFILLER_26_1470 VDD VSS sg13g2f_FILL8
XFILLER_26_1478 VDD VSS sg13g2f_FILL4
XFILLER_26_1496 VDD VSS sg13g2f_FILL2
XFILLER_26_1547 VDD VSS sg13g2f_FILL4
XFILLER_27_430 AVDD VSS sg13g2f_FILL4
XFILLER_27_498 AVDD VSS sg13g2f_FILL8
XFILLER_27_506 AVDD VSS sg13g2f_FILL2
XFILLER_27_513 AVDD VSS sg13g2f_FILL4
XFILLER_27_613 AVDD VSS sg13g2f_FILL8
XFILLER_27_621 AVDD VSS sg13g2f_FILL8
XFILLER_27_629 AVDD VSS sg13g2f_FILL2
XFILLER_27_631 AVDD VSS sg13g2f_FILL1
XFILLER_27_665 AVDD VSS sg13g2f_FILL1
XFILLER_27_746 AVDD VSS sg13g2f_FILL8
XFILLER_27_754 AVDD VSS sg13g2f_FILL2
XFILLER_27_831 AVDD VSS sg13g2f_FILL4
XFILLER_27_835 AVDD VSS sg13g2f_FILL2
XFILLER_27_860 AVDD VSS sg13g2f_FILL8
XFILLER_27_868 AVDD VSS sg13g2f_FILL8
XFILLER_27_876 AVDD VSS sg13g2f_FILL4
XFILLER_27_880 AVDD VSS sg13g2f_FILL2
XFILLER_27_907 AVDD VSS sg13g2f_FILL8
XFILLER_27_915 AVDD VSS sg13g2f_FILL2
XFILLER_27_917 AVDD VSS sg13g2f_FILL1
XFILLER_27_987 AVDD VSS sg13g2f_FILL8
XFILLER_27_995 AVDD VSS sg13g2f_FILL8
XFILLER_27_1003 AVDD VSS sg13g2f_FILL4
XFILLER_27_1007 AVDD VSS sg13g2f_FILL2
XFILLER_27_1020 AVDD VSS sg13g2f_FILL2
XFILLER_27_1022 AVDD VSS sg13g2f_FILL1
XFILLER_27_1066 AVDD VSS sg13g2f_FILL2
XFILLER_27_1118 AVDD VSS sg13g2f_FILL8
XFILLER_27_1126 AVDD VSS sg13g2f_FILL2
XFILLER_27_1192 AVDD VSS sg13g2f_FILL8
XFILLER_27_1200 AVDD VSS sg13g2f_FILL8
XFILLER_27_1208 AVDD VSS sg13g2f_FILL8
XFILLER_27_1216 AVDD VSS sg13g2f_FILL8
XFILLER_27_1224 AVDD VSS sg13g2f_FILL8
XFILLER_27_1232 AVDD VSS sg13g2f_FILL8
XFILLER_27_1240 AVDD VSS sg13g2f_FILL8
XFILLER_27_1248 AVDD VSS sg13g2f_FILL8
XFILLER_27_1256 AVDD VSS sg13g2f_FILL8
XFILLER_27_1264 AVDD VSS sg13g2f_FILL4
XFILLER_27_1390 VDD VSS sg13g2f_FILL8
XFILLER_27_1398 VDD VSS sg13g2f_FILL8
XFILLER_27_1406 VDD VSS sg13g2f_FILL8
XFILLER_27_1414 VDD VSS sg13g2f_FILL8
XFILLER_27_1422 VDD VSS sg13g2f_FILL8
XFILLER_27_1430 VDD VSS sg13g2f_FILL8
XFILLER_27_1438 VDD VSS sg13g2f_FILL8
XFILLER_27_1446 VDD VSS sg13g2f_FILL8
XFILLER_27_1454 VDD VSS sg13g2f_FILL8
XFILLER_27_1462 VDD VSS sg13g2f_FILL8
XFILLER_27_1470 VDD VSS sg13g2f_FILL4
XFILLER_27_1516 VDD VSS sg13g2f_FILL8
XFILLER_27_1524 VDD VSS sg13g2f_FILL8
XFILLER_27_1532 VDD VSS sg13g2f_FILL8
XFILLER_27_1540 VDD VSS sg13g2f_FILL8
XFILLER_27_1548 VDD VSS sg13g2f_FILL2
XFILLER_27_1550 VDD VSS sg13g2f_FILL1
XFILLER_28_7 AVDD VSS sg13g2f_FILL4
XFILLER_28_11 AVDD VSS sg13g2f_FILL2
XFILLER_28_124 AVDD VSS sg13g2f_FILL8
XFILLER_28_132 AVDD VSS sg13g2f_FILL4
XFILLER_28_136 AVDD VSS sg13g2f_FILL2
XFILLER_28_138 AVDD VSS sg13g2f_FILL1
XFILLER_28_155 AVDD VSS sg13g2f_FILL2
XFILLER_28_190 AVDD VSS sg13g2f_FILL8
XFILLER_28_198 AVDD VSS sg13g2f_FILL8
XFILLER_28_206 AVDD VSS sg13g2f_FILL8
XFILLER_28_214 AVDD VSS sg13g2f_FILL8
XFILLER_28_222 AVDD VSS sg13g2f_FILL2
XFILLER_28_231 AVDD VSS sg13g2f_FILL8
XFILLER_28_239 AVDD VSS sg13g2f_FILL8
XFILLER_28_247 AVDD VSS sg13g2f_FILL8
XFILLER_28_255 AVDD VSS sg13g2f_FILL8
XFILLER_28_263 AVDD VSS sg13g2f_FILL8
XFILLER_28_271 AVDD VSS sg13g2f_FILL8
XFILLER_28_279 AVDD VSS sg13g2f_FILL8
XFILLER_28_287 AVDD VSS sg13g2f_FILL4
XFILLER_28_291 AVDD VSS sg13g2f_FILL2
XFILLER_28_293 AVDD VSS sg13g2f_FILL1
XFILLER_28_305 AVDD VSS sg13g2f_FILL8
XFILLER_28_313 AVDD VSS sg13g2f_FILL8
XFILLER_28_321 AVDD VSS sg13g2f_FILL8
XFILLER_28_329 AVDD VSS sg13g2f_FILL4
XFILLER_28_333 AVDD VSS sg13g2f_FILL2
XFILLER_28_335 AVDD VSS sg13g2f_FILL1
XFILLER_28_343 AVDD VSS sg13g2f_FILL4
XFILLER_28_374 AVDD VSS sg13g2f_FILL8
XFILLER_28_382 AVDD VSS sg13g2f_FILL2
XFILLER_28_455 AVDD VSS sg13g2f_FILL8
XFILLER_28_463 AVDD VSS sg13g2f_FILL1
XFILLER_28_496 AVDD VSS sg13g2f_FILL8
XFILLER_28_504 AVDD VSS sg13g2f_FILL8
XFILLER_28_512 AVDD VSS sg13g2f_FILL8
XFILLER_28_520 AVDD VSS sg13g2f_FILL4
XFILLER_28_567 AVDD VSS sg13g2f_FILL4
XFILLER_28_571 AVDD VSS sg13g2f_FILL2
XFILLER_28_573 AVDD VSS sg13g2f_FILL1
XFILLER_28_593 AVDD VSS sg13g2f_FILL4
XFILLER_28_597 AVDD VSS sg13g2f_FILL1
XFILLER_28_617 AVDD VSS sg13g2f_FILL8
XFILLER_28_625 AVDD VSS sg13g2f_FILL4
XFILLER_28_629 AVDD VSS sg13g2f_FILL2
XFILLER_28_631 AVDD VSS sg13g2f_FILL1
XFILLER_28_643 AVDD VSS sg13g2f_FILL8
XFILLER_28_651 AVDD VSS sg13g2f_FILL2
XFILLER_28_653 AVDD VSS sg13g2f_FILL1
XFILLER_28_670 AVDD VSS sg13g2f_FILL2
XFILLER_28_743 AVDD VSS sg13g2f_FILL8
XFILLER_28_751 AVDD VSS sg13g2f_FILL4
XFILLER_28_755 AVDD VSS sg13g2f_FILL1
XFILLER_28_778 AVDD VSS sg13g2f_FILL4
XFILLER_28_782 AVDD VSS sg13g2f_FILL2
XFILLER_28_791 AVDD VSS sg13g2f_FILL8
XFILLER_28_799 AVDD VSS sg13g2f_FILL4
XFILLER_28_803 AVDD VSS sg13g2f_FILL2
XFILLER_28_805 AVDD VSS sg13g2f_FILL1
XFILLER_28_870 AVDD VSS sg13g2f_FILL8
XFILLER_28_878 AVDD VSS sg13g2f_FILL2
XFILLER_28_891 AVDD VSS sg13g2f_FILL4
XFILLER_28_895 AVDD VSS sg13g2f_FILL1
XFILLER_28_914 AVDD VSS sg13g2f_FILL1
XFILLER_28_990 AVDD VSS sg13g2f_FILL8
XFILLER_28_998 AVDD VSS sg13g2f_FILL8
XFILLER_28_1006 AVDD VSS sg13g2f_FILL2
XFILLER_28_1015 AVDD VSS sg13g2f_FILL1
XFILLER_28_1059 AVDD VSS sg13g2f_FILL4
XFILLER_28_1063 AVDD VSS sg13g2f_FILL2
XFILLER_28_1081 AVDD VSS sg13g2f_FILL1
XFILLER_28_1118 AVDD VSS sg13g2f_FILL2
XFILLER_28_1127 AVDD VSS sg13g2f_FILL1
XFILLER_28_1182 AVDD VSS sg13g2f_FILL8
XFILLER_28_1190 AVDD VSS sg13g2f_FILL8
XFILLER_28_1198 AVDD VSS sg13g2f_FILL8
XFILLER_28_1206 AVDD VSS sg13g2f_FILL8
XFILLER_28_1214 AVDD VSS sg13g2f_FILL8
XFILLER_28_1222 AVDD VSS sg13g2f_FILL8
XFILLER_28_1230 AVDD VSS sg13g2f_FILL2
XFILLER_28_1239 AVDD VSS sg13g2f_FILL8
XFILLER_28_1247 AVDD VSS sg13g2f_FILL8
XFILLER_28_1255 AVDD VSS sg13g2f_FILL8
XFILLER_28_1263 AVDD VSS sg13g2f_FILL4
XFILLER_28_1267 AVDD VSS sg13g2f_FILL1
XFILLER_28_1390 VDD VSS sg13g2f_FILL8
XFILLER_28_1398 VDD VSS sg13g2f_FILL8
XFILLER_28_1406 VDD VSS sg13g2f_FILL8
XFILLER_28_1414 VDD VSS sg13g2f_FILL8
XFILLER_28_1422 VDD VSS sg13g2f_FILL8
XFILLER_28_1430 VDD VSS sg13g2f_FILL8
XFILLER_28_1438 VDD VSS sg13g2f_FILL8
XFILLER_28_1446 VDD VSS sg13g2f_FILL8
XFILLER_28_1454 VDD VSS sg13g2f_FILL8
XFILLER_28_1462 VDD VSS sg13g2f_FILL8
XFILLER_28_1470 VDD VSS sg13g2f_FILL8
XFILLER_28_1478 VDD VSS sg13g2f_FILL8
XFILLER_28_1486 VDD VSS sg13g2f_FILL1
XFILLER_28_1513 VDD VSS sg13g2f_FILL8
XFILLER_28_1521 VDD VSS sg13g2f_FILL8
XFILLER_28_1529 VDD VSS sg13g2f_FILL8
XFILLER_28_1537 VDD VSS sg13g2f_FILL8
XFILLER_28_1545 VDD VSS sg13g2f_FILL4
XFILLER_28_1549 VDD VSS sg13g2f_FILL2
XFILLER_29_7 AVDD VSS sg13g2f_FILL4
XFILLER_29_11 AVDD VSS sg13g2f_FILL1
XFILLER_29_76 AVDD VSS sg13g2f_FILL8
XFILLER_29_84 AVDD VSS sg13g2f_FILL8
XFILLER_29_92 AVDD VSS sg13g2f_FILL8
XFILLER_29_100 AVDD VSS sg13g2f_FILL8
XFILLER_29_108 AVDD VSS sg13g2f_FILL8
XFILLER_29_116 AVDD VSS sg13g2f_FILL8
XFILLER_29_124 AVDD VSS sg13g2f_FILL8
XFILLER_29_132 AVDD VSS sg13g2f_FILL4
XFILLER_29_152 AVDD VSS sg13g2f_FILL4
XFILLER_29_156 AVDD VSS sg13g2f_FILL1
XFILLER_29_168 AVDD VSS sg13g2f_FILL8
XFILLER_29_176 AVDD VSS sg13g2f_FILL8
XFILLER_29_184 AVDD VSS sg13g2f_FILL8
XFILLER_29_192 AVDD VSS sg13g2f_FILL8
XFILLER_29_200 AVDD VSS sg13g2f_FILL8
XFILLER_29_208 AVDD VSS sg13g2f_FILL8
XFILLER_29_216 AVDD VSS sg13g2f_FILL8
XFILLER_29_224 AVDD VSS sg13g2f_FILL4
XFILLER_29_228 AVDD VSS sg13g2f_FILL2
XFILLER_29_230 AVDD VSS sg13g2f_FILL1
XFILLER_29_238 AVDD VSS sg13g2f_FILL8
XFILLER_29_246 AVDD VSS sg13g2f_FILL8
XFILLER_29_254 AVDD VSS sg13g2f_FILL8
XFILLER_29_262 AVDD VSS sg13g2f_FILL8
XFILLER_29_270 AVDD VSS sg13g2f_FILL8
XFILLER_29_278 AVDD VSS sg13g2f_FILL8
XFILLER_29_286 AVDD VSS sg13g2f_FILL8
XFILLER_29_294 AVDD VSS sg13g2f_FILL8
XFILLER_29_302 AVDD VSS sg13g2f_FILL8
XFILLER_29_310 AVDD VSS sg13g2f_FILL8
XFILLER_29_318 AVDD VSS sg13g2f_FILL8
XFILLER_29_326 AVDD VSS sg13g2f_FILL8
XFILLER_29_334 AVDD VSS sg13g2f_FILL8
XFILLER_29_342 AVDD VSS sg13g2f_FILL8
XFILLER_29_350 AVDD VSS sg13g2f_FILL8
XFILLER_29_358 AVDD VSS sg13g2f_FILL1
XFILLER_29_364 AVDD VSS sg13g2f_FILL8
XFILLER_29_372 AVDD VSS sg13g2f_FILL8
XFILLER_29_380 AVDD VSS sg13g2f_FILL4
XFILLER_29_448 AVDD VSS sg13g2f_FILL2
XFILLER_29_450 AVDD VSS sg13g2f_FILL1
XFILLER_29_485 AVDD VSS sg13g2f_FILL8
XFILLER_29_493 AVDD VSS sg13g2f_FILL8
XFILLER_29_501 AVDD VSS sg13g2f_FILL8
XFILLER_29_509 AVDD VSS sg13g2f_FILL4
XFILLER_29_593 AVDD VSS sg13g2f_FILL4
XFILLER_29_613 AVDD VSS sg13g2f_FILL8
XFILLER_29_621 AVDD VSS sg13g2f_FILL8
XFILLER_29_629 AVDD VSS sg13g2f_FILL8
XFILLER_29_637 AVDD VSS sg13g2f_FILL8
XFILLER_29_645 AVDD VSS sg13g2f_FILL8
XFILLER_29_653 AVDD VSS sg13g2f_FILL8
XFILLER_29_661 AVDD VSS sg13g2f_FILL1
XFILLER_29_673 AVDD VSS sg13g2f_FILL4
XFILLER_29_741 AVDD VSS sg13g2f_FILL8
XFILLER_29_749 AVDD VSS sg13g2f_FILL8
XFILLER_29_757 AVDD VSS sg13g2f_FILL8
XFILLER_29_765 AVDD VSS sg13g2f_FILL8
XFILLER_29_773 AVDD VSS sg13g2f_FILL8
XFILLER_29_781 AVDD VSS sg13g2f_FILL8
XFILLER_29_789 AVDD VSS sg13g2f_FILL4
XFILLER_29_793 AVDD VSS sg13g2f_FILL2
XFILLER_29_827 AVDD VSS sg13g2f_FILL2
XFILLER_29_829 AVDD VSS sg13g2f_FILL1
XFILLER_29_855 AVDD VSS sg13g2f_FILL2
XFILLER_29_868 AVDD VSS sg13g2f_FILL8
XFILLER_29_876 AVDD VSS sg13g2f_FILL8
XFILLER_29_909 AVDD VSS sg13g2f_FILL4
XFILLER_29_931 AVDD VSS sg13g2f_FILL8
XFILLER_29_939 AVDD VSS sg13g2f_FILL8
XFILLER_29_947 AVDD VSS sg13g2f_FILL1
XFILLER_29_991 AVDD VSS sg13g2f_FILL8
XFILLER_29_999 AVDD VSS sg13g2f_FILL8
XFILLER_29_1007 AVDD VSS sg13g2f_FILL4
XFILLER_29_1011 AVDD VSS sg13g2f_FILL2
XFILLER_29_1013 AVDD VSS sg13g2f_FILL1
XFILLER_29_1047 AVDD VSS sg13g2f_FILL8
XFILLER_29_1055 AVDD VSS sg13g2f_FILL8
XFILLER_29_1063 AVDD VSS sg13g2f_FILL8
XFILLER_29_1071 AVDD VSS sg13g2f_FILL4
XFILLER_29_1118 AVDD VSS sg13g2f_FILL8
XFILLER_29_1126 AVDD VSS sg13g2f_FILL8
XFILLER_29_1134 AVDD VSS sg13g2f_FILL1
XFILLER_29_1151 AVDD VSS sg13g2f_FILL4
XFILLER_29_1173 AVDD VSS sg13g2f_FILL8
XFILLER_29_1181 AVDD VSS sg13g2f_FILL8
XFILLER_29_1189 AVDD VSS sg13g2f_FILL8
XFILLER_29_1197 AVDD VSS sg13g2f_FILL8
XFILLER_29_1205 AVDD VSS sg13g2f_FILL8
XFILLER_29_1213 AVDD VSS sg13g2f_FILL8
XFILLER_29_1221 AVDD VSS sg13g2f_FILL8
XFILLER_29_1229 AVDD VSS sg13g2f_FILL8
XFILLER_29_1237 AVDD VSS sg13g2f_FILL8
XFILLER_29_1245 AVDD VSS sg13g2f_FILL8
XFILLER_29_1253 AVDD VSS sg13g2f_FILL8
XFILLER_29_1261 AVDD VSS sg13g2f_FILL4
XFILLER_29_1265 AVDD VSS sg13g2f_FILL2
XFILLER_29_1267 AVDD VSS sg13g2f_FILL1
XFILLER_29_1390 VDD VSS sg13g2f_FILL8
XFILLER_29_1398 VDD VSS sg13g2f_FILL8
XFILLER_29_1406 VDD VSS sg13g2f_FILL8
XFILLER_29_1414 VDD VSS sg13g2f_FILL8
XFILLER_29_1422 VDD VSS sg13g2f_FILL8
XFILLER_29_1430 VDD VSS sg13g2f_FILL8
XFILLER_29_1438 VDD VSS sg13g2f_FILL8
XFILLER_29_1446 VDD VSS sg13g2f_FILL8
XFILLER_29_1454 VDD VSS sg13g2f_FILL8
XFILLER_29_1462 VDD VSS sg13g2f_FILL8
XFILLER_29_1470 VDD VSS sg13g2f_FILL4
XFILLER_29_1474 VDD VSS sg13g2f_FILL1
XFILLER_29_1528 VDD VSS sg13g2f_FILL8
XFILLER_29_1536 VDD VSS sg13g2f_FILL8
XFILLER_29_1544 VDD VSS sg13g2f_FILL4
XFILLER_29_1548 VDD VSS sg13g2f_FILL2
XFILLER_29_1550 VDD VSS sg13g2f_FILL1
XFILLER_30_7 AVDD VSS sg13g2f_FILL8
XFILLER_30_15 AVDD VSS sg13g2f_FILL8
XFILLER_30_23 AVDD VSS sg13g2f_FILL2
XFILLER_30_25 AVDD VSS sg13g2f_FILL1
XFILLER_30_47 AVDD VSS sg13g2f_FILL1
XFILLER_30_119 AVDD VSS sg13g2f_FILL8
XFILLER_30_127 AVDD VSS sg13g2f_FILL8
XFILLER_30_135 AVDD VSS sg13g2f_FILL8
XFILLER_30_143 AVDD VSS sg13g2f_FILL8
XFILLER_30_151 AVDD VSS sg13g2f_FILL8
XFILLER_30_159 AVDD VSS sg13g2f_FILL8
XFILLER_30_167 AVDD VSS sg13g2f_FILL8
XFILLER_30_175 AVDD VSS sg13g2f_FILL8
XFILLER_30_183 AVDD VSS sg13g2f_FILL8
XFILLER_30_191 AVDD VSS sg13g2f_FILL8
XFILLER_30_199 AVDD VSS sg13g2f_FILL8
XFILLER_30_207 AVDD VSS sg13g2f_FILL8
XFILLER_30_215 AVDD VSS sg13g2f_FILL8
XFILLER_30_223 AVDD VSS sg13g2f_FILL1
XFILLER_30_231 AVDD VSS sg13g2f_FILL8
XFILLER_30_239 AVDD VSS sg13g2f_FILL8
XFILLER_30_247 AVDD VSS sg13g2f_FILL8
XFILLER_30_255 AVDD VSS sg13g2f_FILL8
XFILLER_30_263 AVDD VSS sg13g2f_FILL8
XFILLER_30_271 AVDD VSS sg13g2f_FILL8
XFILLER_30_279 AVDD VSS sg13g2f_FILL8
XFILLER_30_287 AVDD VSS sg13g2f_FILL8
XFILLER_30_295 AVDD VSS sg13g2f_FILL8
XFILLER_30_303 AVDD VSS sg13g2f_FILL8
XFILLER_30_311 AVDD VSS sg13g2f_FILL8
XFILLER_30_319 AVDD VSS sg13g2f_FILL8
XFILLER_30_327 AVDD VSS sg13g2f_FILL8
XFILLER_30_335 AVDD VSS sg13g2f_FILL1
XFILLER_30_343 AVDD VSS sg13g2f_FILL8
XFILLER_30_351 AVDD VSS sg13g2f_FILL8
XFILLER_30_359 AVDD VSS sg13g2f_FILL8
XFILLER_30_367 AVDD VSS sg13g2f_FILL8
XFILLER_30_375 AVDD VSS sg13g2f_FILL8
XFILLER_30_383 AVDD VSS sg13g2f_FILL1
XFILLER_30_455 AVDD VSS sg13g2f_FILL1
XFILLER_30_467 AVDD VSS sg13g2f_FILL8
XFILLER_30_475 AVDD VSS sg13g2f_FILL8
XFILLER_30_483 AVDD VSS sg13g2f_FILL8
XFILLER_30_491 AVDD VSS sg13g2f_FILL8
XFILLER_30_499 AVDD VSS sg13g2f_FILL8
XFILLER_30_507 AVDD VSS sg13g2f_FILL8
XFILLER_30_515 AVDD VSS sg13g2f_FILL8
XFILLER_30_523 AVDD VSS sg13g2f_FILL8
XFILLER_30_531 AVDD VSS sg13g2f_FILL8
XFILLER_30_539 AVDD VSS sg13g2f_FILL8
XFILLER_30_547 AVDD VSS sg13g2f_FILL8
XFILLER_30_555 AVDD VSS sg13g2f_FILL4
XFILLER_30_559 AVDD VSS sg13g2f_FILL1
XFILLER_30_567 AVDD VSS sg13g2f_FILL8
XFILLER_30_575 AVDD VSS sg13g2f_FILL8
XFILLER_30_583 AVDD VSS sg13g2f_FILL8
XFILLER_30_591 AVDD VSS sg13g2f_FILL8
XFILLER_30_599 AVDD VSS sg13g2f_FILL8
XFILLER_30_607 AVDD VSS sg13g2f_FILL8
XFILLER_30_615 AVDD VSS sg13g2f_FILL8
XFILLER_30_623 AVDD VSS sg13g2f_FILL8
XFILLER_30_631 AVDD VSS sg13g2f_FILL8
XFILLER_30_639 AVDD VSS sg13g2f_FILL8
XFILLER_30_647 AVDD VSS sg13g2f_FILL8
XFILLER_30_655 AVDD VSS sg13g2f_FILL8
XFILLER_30_663 AVDD VSS sg13g2f_FILL8
XFILLER_30_671 AVDD VSS sg13g2f_FILL1
XFILLER_30_679 AVDD VSS sg13g2f_FILL8
XFILLER_30_687 AVDD VSS sg13g2f_FILL8
XFILLER_30_695 AVDD VSS sg13g2f_FILL8
XFILLER_30_714 AVDD VSS sg13g2f_FILL8
XFILLER_30_722 AVDD VSS sg13g2f_FILL8
XFILLER_30_730 AVDD VSS sg13g2f_FILL8
XFILLER_30_738 AVDD VSS sg13g2f_FILL8
XFILLER_30_746 AVDD VSS sg13g2f_FILL8
XFILLER_30_754 AVDD VSS sg13g2f_FILL8
XFILLER_30_762 AVDD VSS sg13g2f_FILL8
XFILLER_30_770 AVDD VSS sg13g2f_FILL8
XFILLER_30_778 AVDD VSS sg13g2f_FILL4
XFILLER_30_782 AVDD VSS sg13g2f_FILL2
XFILLER_30_791 AVDD VSS sg13g2f_FILL8
XFILLER_30_799 AVDD VSS sg13g2f_FILL8
XFILLER_30_807 AVDD VSS sg13g2f_FILL8
XFILLER_30_815 AVDD VSS sg13g2f_FILL8
XFILLER_30_823 AVDD VSS sg13g2f_FILL8
XFILLER_30_831 AVDD VSS sg13g2f_FILL8
XFILLER_30_839 AVDD VSS sg13g2f_FILL8
XFILLER_30_847 AVDD VSS sg13g2f_FILL8
XFILLER_30_855 AVDD VSS sg13g2f_FILL8
XFILLER_30_863 AVDD VSS sg13g2f_FILL8
XFILLER_30_871 AVDD VSS sg13g2f_FILL8
XFILLER_30_879 AVDD VSS sg13g2f_FILL8
XFILLER_30_887 AVDD VSS sg13g2f_FILL8
XFILLER_30_895 AVDD VSS sg13g2f_FILL1
XFILLER_30_903 AVDD VSS sg13g2f_FILL8
XFILLER_30_911 AVDD VSS sg13g2f_FILL8
XFILLER_30_919 AVDD VSS sg13g2f_FILL8
XFILLER_30_927 AVDD VSS sg13g2f_FILL8
XFILLER_30_935 AVDD VSS sg13g2f_FILL8
XFILLER_30_943 AVDD VSS sg13g2f_FILL8
XFILLER_30_951 AVDD VSS sg13g2f_FILL8
XFILLER_30_959 AVDD VSS sg13g2f_FILL8
XFILLER_30_967 AVDD VSS sg13g2f_FILL1
XFILLER_30_979 AVDD VSS sg13g2f_FILL8
XFILLER_30_987 AVDD VSS sg13g2f_FILL8
XFILLER_30_995 AVDD VSS sg13g2f_FILL8
XFILLER_30_1003 AVDD VSS sg13g2f_FILL4
XFILLER_30_1007 AVDD VSS sg13g2f_FILL1
XFILLER_30_1015 AVDD VSS sg13g2f_FILL8
XFILLER_30_1023 AVDD VSS sg13g2f_FILL8
XFILLER_30_1031 AVDD VSS sg13g2f_FILL8
XFILLER_30_1039 AVDD VSS sg13g2f_FILL8
XFILLER_30_1047 AVDD VSS sg13g2f_FILL8
XFILLER_30_1055 AVDD VSS sg13g2f_FILL8
XFILLER_30_1063 AVDD VSS sg13g2f_FILL8
XFILLER_30_1071 AVDD VSS sg13g2f_FILL8
XFILLER_30_1079 AVDD VSS sg13g2f_FILL8
XFILLER_30_1087 AVDD VSS sg13g2f_FILL8
XFILLER_30_1095 AVDD VSS sg13g2f_FILL8
XFILLER_30_1103 AVDD VSS sg13g2f_FILL8
XFILLER_30_1111 AVDD VSS sg13g2f_FILL8
XFILLER_30_1119 AVDD VSS sg13g2f_FILL1
XFILLER_30_1127 AVDD VSS sg13g2f_FILL8
XFILLER_30_1135 AVDD VSS sg13g2f_FILL8
XFILLER_30_1143 AVDD VSS sg13g2f_FILL8
XFILLER_30_1151 AVDD VSS sg13g2f_FILL8
XFILLER_30_1159 AVDD VSS sg13g2f_FILL8
XFILLER_30_1167 AVDD VSS sg13g2f_FILL8
XFILLER_30_1175 AVDD VSS sg13g2f_FILL8
XFILLER_30_1183 AVDD VSS sg13g2f_FILL8
XFILLER_30_1191 AVDD VSS sg13g2f_FILL8
XFILLER_30_1199 AVDD VSS sg13g2f_FILL8
XFILLER_30_1207 AVDD VSS sg13g2f_FILL8
XFILLER_30_1215 AVDD VSS sg13g2f_FILL8
XFILLER_30_1223 AVDD VSS sg13g2f_FILL8
XFILLER_30_1231 AVDD VSS sg13g2f_FILL1
XFILLER_30_1239 AVDD VSS sg13g2f_FILL8
XFILLER_30_1247 AVDD VSS sg13g2f_FILL8
XFILLER_30_1255 AVDD VSS sg13g2f_FILL8
XFILLER_30_1263 AVDD VSS sg13g2f_FILL4
XFILLER_30_1267 AVDD VSS sg13g2f_FILL1
XFILLER_30_1390 VDD VSS sg13g2f_FILL8
XFILLER_30_1398 VDD VSS sg13g2f_FILL8
XFILLER_30_1406 VDD VSS sg13g2f_FILL8
XFILLER_30_1414 VDD VSS sg13g2f_FILL8
XFILLER_30_1422 VDD VSS sg13g2f_FILL8
XFILLER_30_1430 VDD VSS sg13g2f_FILL8
XFILLER_30_1438 VDD VSS sg13g2f_FILL8
XFILLER_30_1446 VDD VSS sg13g2f_FILL8
XFILLER_30_1454 VDD VSS sg13g2f_FILL2
XFILLER_30_1547 VDD VSS sg13g2f_FILL4
XFILLER_31_1390 VDD VSS sg13g2f_FILL8
XFILLER_31_1398 VDD VSS sg13g2f_FILL8
XFILLER_31_1406 VDD VSS sg13g2f_FILL8
XFILLER_31_1414 VDD VSS sg13g2f_FILL8
XFILLER_31_1422 VDD VSS sg13g2f_FILL8
XFILLER_31_1430 VDD VSS sg13g2f_FILL8
XFILLER_31_1438 VDD VSS sg13g2f_FILL8
XFILLER_31_1446 VDD VSS sg13g2f_FILL8
XFILLER_31_1454 VDD VSS sg13g2f_FILL8
XFILLER_31_1462 VDD VSS sg13g2f_FILL8
XFILLER_31_1470 VDD VSS sg13g2f_FILL8
XFILLER_31_1478 VDD VSS sg13g2f_FILL8
XFILLER_31_1486 VDD VSS sg13g2f_FILL8
XFILLER_31_1494 VDD VSS sg13g2f_FILL8
XFILLER_31_1502 VDD VSS sg13g2f_FILL4
XFILLER_31_1517 VDD VSS sg13g2f_FILL8
XFILLER_31_1525 VDD VSS sg13g2f_FILL8
XFILLER_31_1533 VDD VSS sg13g2f_FILL8
XFILLER_31_1541 VDD VSS sg13g2f_FILL8
XFILLER_31_1549 VDD VSS sg13g2f_FILL2
XFILLER_32_1390 VDD VSS sg13g2f_FILL8
XFILLER_32_1398 VDD VSS sg13g2f_FILL8
XFILLER_32_1406 VDD VSS sg13g2f_FILL8
XFILLER_32_1414 VDD VSS sg13g2f_FILL8
XFILLER_32_1422 VDD VSS sg13g2f_FILL8
XFILLER_32_1430 VDD VSS sg13g2f_FILL8
XFILLER_32_1438 VDD VSS sg13g2f_FILL8
XFILLER_32_1446 VDD VSS sg13g2f_FILL8
XFILLER_32_1454 VDD VSS sg13g2f_FILL8
XFILLER_32_1462 VDD VSS sg13g2f_FILL8
XFILLER_32_1470 VDD VSS sg13g2f_FILL8
XFILLER_32_1478 VDD VSS sg13g2f_FILL8
XFILLER_32_1486 VDD VSS sg13g2f_FILL8
XFILLER_32_1494 VDD VSS sg13g2f_FILL4
XFILLER_32_1516 VDD VSS sg13g2f_FILL8
XFILLER_32_1524 VDD VSS sg13g2f_FILL8
XFILLER_32_1532 VDD VSS sg13g2f_FILL8
XFILLER_32_1540 VDD VSS sg13g2f_FILL8
XFILLER_32_1548 VDD VSS sg13g2f_FILL2
XFILLER_32_1550 VDD VSS sg13g2f_FILL1
XFILLER_33_1390 VDD VSS sg13g2f_FILL8
XFILLER_33_1398 VDD VSS sg13g2f_FILL8
XFILLER_33_1406 VDD VSS sg13g2f_FILL8
XFILLER_33_1414 VDD VSS sg13g2f_FILL8
XFILLER_33_1422 VDD VSS sg13g2f_FILL8
XFILLER_33_1430 VDD VSS sg13g2f_FILL8
XFILLER_33_1438 VDD VSS sg13g2f_FILL8
XFILLER_33_1446 VDD VSS sg13g2f_FILL8
XFILLER_33_1454 VDD VSS sg13g2f_FILL8
XFILLER_33_1462 VDD VSS sg13g2f_FILL8
XFILLER_33_1470 VDD VSS sg13g2f_FILL4
XFILLER_33_1474 VDD VSS sg13g2f_FILL1
XFILLER_33_1531 VDD VSS sg13g2f_FILL8
XFILLER_33_1539 VDD VSS sg13g2f_FILL8
XFILLER_33_1547 VDD VSS sg13g2f_FILL4
XFILLER_34_1390 VDD VSS sg13g2f_FILL8
XFILLER_34_1398 VDD VSS sg13g2f_FILL8
XFILLER_34_1406 VDD VSS sg13g2f_FILL8
XFILLER_34_1414 VDD VSS sg13g2f_FILL8
XFILLER_34_1422 VDD VSS sg13g2f_FILL8
XFILLER_34_1430 VDD VSS sg13g2f_FILL8
XFILLER_34_1438 VDD VSS sg13g2f_FILL8
XFILLER_34_1446 VDD VSS sg13g2f_FILL8
XFILLER_34_1454 VDD VSS sg13g2f_FILL8
XFILLER_34_1462 VDD VSS sg13g2f_FILL8
XFILLER_34_1470 VDD VSS sg13g2f_FILL8
XFILLER_34_1478 VDD VSS sg13g2f_FILL8
XFILLER_34_1486 VDD VSS sg13g2f_FILL8
XFILLER_34_1494 VDD VSS sg13g2f_FILL4
XFILLER_34_1505 VDD VSS sg13g2f_FILL4
XFILLER_34_1520 VDD VSS sg13g2f_FILL8
XFILLER_34_1528 VDD VSS sg13g2f_FILL8
XFILLER_34_1536 VDD VSS sg13g2f_FILL8
XFILLER_34_1544 VDD VSS sg13g2f_FILL4
XFILLER_34_1548 VDD VSS sg13g2f_FILL2
XFILLER_34_1550 VDD VSS sg13g2f_FILL1
XFILLER_35_1390 VDD VSS sg13g2f_FILL8
XFILLER_35_1398 VDD VSS sg13g2f_FILL8
XFILLER_35_1406 VDD VSS sg13g2f_FILL8
XFILLER_35_1414 VDD VSS sg13g2f_FILL8
XFILLER_35_1422 VDD VSS sg13g2f_FILL8
XFILLER_35_1430 VDD VSS sg13g2f_FILL8
XFILLER_35_1438 VDD VSS sg13g2f_FILL8
XFILLER_35_1446 VDD VSS sg13g2f_FILL8
XFILLER_35_1454 VDD VSS sg13g2f_FILL8
XFILLER_35_1462 VDD VSS sg13g2f_FILL8
XFILLER_35_1470 VDD VSS sg13g2f_FILL8
XFILLER_35_1478 VDD VSS sg13g2f_FILL8
XFILLER_35_1486 VDD VSS sg13g2f_FILL8
XFILLER_35_1536 VDD VSS sg13g2f_FILL8
XFILLER_35_1544 VDD VSS sg13g2f_FILL4
XFILLER_35_1548 VDD VSS sg13g2f_FILL2
XFILLER_35_1550 VDD VSS sg13g2f_FILL1
XFILLER_36_1390 VDD VSS sg13g2f_FILL8
XFILLER_36_1398 VDD VSS sg13g2f_FILL8
XFILLER_36_1406 VDD VSS sg13g2f_FILL8
XFILLER_36_1414 VDD VSS sg13g2f_FILL8
XFILLER_36_1422 VDD VSS sg13g2f_FILL8
XFILLER_36_1430 VDD VSS sg13g2f_FILL8
XFILLER_36_1438 VDD VSS sg13g2f_FILL8
XFILLER_36_1446 VDD VSS sg13g2f_FILL8
XFILLER_36_1454 VDD VSS sg13g2f_FILL8
XFILLER_36_1462 VDD VSS sg13g2f_FILL8
XFILLER_36_1470 VDD VSS sg13g2f_FILL8
XFILLER_36_1478 VDD VSS sg13g2f_FILL8
XFILLER_36_1486 VDD VSS sg13g2f_FILL8
XFILLER_36_1494 VDD VSS sg13g2f_FILL4
XFILLER_36_1505 VDD VSS sg13g2f_FILL4
XFILLER_36_1509 VDD VSS sg13g2f_FILL2
XFILLER_36_1511 VDD VSS sg13g2f_FILL1
XFILLER_36_1545 VDD VSS sg13g2f_FILL4
XFILLER_36_1549 VDD VSS sg13g2f_FILL2
XFILLER_37_1390 VDD VSS sg13g2f_FILL8
XFILLER_37_1398 VDD VSS sg13g2f_FILL8
XFILLER_37_1406 VDD VSS sg13g2f_FILL8
XFILLER_37_1414 VDD VSS sg13g2f_FILL8
XFILLER_37_1422 VDD VSS sg13g2f_FILL8
XFILLER_37_1430 VDD VSS sg13g2f_FILL8
XFILLER_37_1438 VDD VSS sg13g2f_FILL8
XFILLER_37_1446 VDD VSS sg13g2f_FILL8
XFILLER_37_1454 VDD VSS sg13g2f_FILL8
XFILLER_37_1462 VDD VSS sg13g2f_FILL8
XFILLER_37_1470 VDD VSS sg13g2f_FILL8
XFILLER_37_1478 VDD VSS sg13g2f_FILL8
XFILLER_37_1486 VDD VSS sg13g2f_FILL8
XFILLER_37_1494 VDD VSS sg13g2f_FILL8
XFILLER_37_1502 VDD VSS sg13g2f_FILL8
XFILLER_37_1510 VDD VSS sg13g2f_FILL4
XFILLER_37_1525 VDD VSS sg13g2f_FILL8
XFILLER_37_1533 VDD VSS sg13g2f_FILL8
XFILLER_37_1541 VDD VSS sg13g2f_FILL8
XFILLER_37_1549 VDD VSS sg13g2f_FILL2
XFILLER_38_1390 VDD VSS sg13g2f_FILL8
XFILLER_38_1398 VDD VSS sg13g2f_FILL8
XFILLER_38_1406 VDD VSS sg13g2f_FILL8
XFILLER_38_1414 VDD VSS sg13g2f_FILL8
XFILLER_38_1422 VDD VSS sg13g2f_FILL8
XFILLER_38_1430 VDD VSS sg13g2f_FILL8
XFILLER_38_1438 VDD VSS sg13g2f_FILL8
XFILLER_38_1446 VDD VSS sg13g2f_FILL8
XFILLER_38_1454 VDD VSS sg13g2f_FILL8
XFILLER_38_1462 VDD VSS sg13g2f_FILL8
XFILLER_38_1470 VDD VSS sg13g2f_FILL8
XFILLER_38_1478 VDD VSS sg13g2f_FILL8
XFILLER_38_1486 VDD VSS sg13g2f_FILL8
XFILLER_38_1494 VDD VSS sg13g2f_FILL4
XFILLER_38_1505 VDD VSS sg13g2f_FILL8
XFILLER_38_1513 VDD VSS sg13g2f_FILL1
XFILLER_38_1528 VDD VSS sg13g2f_FILL8
XFILLER_38_1536 VDD VSS sg13g2f_FILL8
XFILLER_38_1544 VDD VSS sg13g2f_FILL4
XFILLER_38_1548 VDD VSS sg13g2f_FILL2
XFILLER_38_1550 VDD VSS sg13g2f_FILL1
XFILLER_39_1390 VDD VSS sg13g2f_FILL8
XFILLER_39_1398 VDD VSS sg13g2f_FILL8
XFILLER_39_1406 VDD VSS sg13g2f_FILL8
XFILLER_39_1414 VDD VSS sg13g2f_FILL8
XFILLER_39_1422 VDD VSS sg13g2f_FILL8
XFILLER_39_1430 VDD VSS sg13g2f_FILL8
XFILLER_39_1438 VDD VSS sg13g2f_FILL8
XFILLER_39_1446 VDD VSS sg13g2f_FILL8
XFILLER_39_1454 VDD VSS sg13g2f_FILL8
XFILLER_39_1462 VDD VSS sg13g2f_FILL8
XFILLER_39_1470 VDD VSS sg13g2f_FILL8
XFILLER_39_1478 VDD VSS sg13g2f_FILL8
XFILLER_39_1486 VDD VSS sg13g2f_FILL8
XFILLER_39_1494 VDD VSS sg13g2f_FILL8
XFILLER_39_1502 VDD VSS sg13g2f_FILL8
XFILLER_39_1510 VDD VSS sg13g2f_FILL4
XFILLER_39_1514 VDD VSS sg13g2f_FILL1
XFILLER_39_1526 VDD VSS sg13g2f_FILL8
XFILLER_39_1534 VDD VSS sg13g2f_FILL8
XFILLER_39_1542 VDD VSS sg13g2f_FILL8
XFILLER_39_1550 VDD VSS sg13g2f_FILL1
XFILLER_40_1390 VDD VSS sg13g2f_FILL8
XFILLER_40_1398 VDD VSS sg13g2f_FILL8
XFILLER_40_1406 VDD VSS sg13g2f_FILL8
XFILLER_40_1414 VDD VSS sg13g2f_FILL8
XFILLER_40_1422 VDD VSS sg13g2f_FILL8
XFILLER_40_1430 VDD VSS sg13g2f_FILL8
XFILLER_40_1438 VDD VSS sg13g2f_FILL8
XFILLER_40_1446 VDD VSS sg13g2f_FILL8
XFILLER_40_1454 VDD VSS sg13g2f_FILL8
XFILLER_40_1462 VDD VSS sg13g2f_FILL8
XFILLER_40_1470 VDD VSS sg13g2f_FILL8
XFILLER_40_1478 VDD VSS sg13g2f_FILL8
XFILLER_40_1486 VDD VSS sg13g2f_FILL8
XFILLER_40_1494 VDD VSS sg13g2f_FILL4
XFILLER_40_1505 VDD VSS sg13g2f_FILL8
XFILLER_40_1513 VDD VSS sg13g2f_FILL4
XFILLER_40_1517 VDD VSS sg13g2f_FILL1
XFILLER_40_1529 VDD VSS sg13g2f_FILL8
XFILLER_40_1537 VDD VSS sg13g2f_FILL8
XFILLER_40_1545 VDD VSS sg13g2f_FILL4
XFILLER_40_1549 VDD VSS sg13g2f_FILL2
XFILLER_41_1390 VDD VSS sg13g2f_FILL8
XFILLER_41_1398 VDD VSS sg13g2f_FILL8
XFILLER_41_1406 VDD VSS sg13g2f_FILL8
XFILLER_41_1414 VDD VSS sg13g2f_FILL8
XFILLER_41_1422 VDD VSS sg13g2f_FILL8
XFILLER_41_1430 VDD VSS sg13g2f_FILL8
XFILLER_41_1438 VDD VSS sg13g2f_FILL8
XFILLER_41_1446 VDD VSS sg13g2f_FILL8
XFILLER_41_1454 VDD VSS sg13g2f_FILL8
XFILLER_41_1462 VDD VSS sg13g2f_FILL8
XFILLER_41_1470 VDD VSS sg13g2f_FILL8
XFILLER_41_1478 VDD VSS sg13g2f_FILL8
XFILLER_41_1486 VDD VSS sg13g2f_FILL8
XFILLER_41_1494 VDD VSS sg13g2f_FILL8
XFILLER_41_1502 VDD VSS sg13g2f_FILL8
XFILLER_41_1510 VDD VSS sg13g2f_FILL2
XFILLER_41_1512 VDD VSS sg13g2f_FILL1
XFILLER_41_1534 VDD VSS sg13g2f_FILL8
XFILLER_41_1542 VDD VSS sg13g2f_FILL8
XFILLER_41_1550 VDD VSS sg13g2f_FILL1
XFILLER_42_1390 VDD VSS sg13g2f_FILL8
XFILLER_42_1398 VDD VSS sg13g2f_FILL8
XFILLER_42_1406 VDD VSS sg13g2f_FILL8
XFILLER_42_1414 VDD VSS sg13g2f_FILL8
XFILLER_42_1422 VDD VSS sg13g2f_FILL8
XFILLER_42_1430 VDD VSS sg13g2f_FILL8
XFILLER_42_1438 VDD VSS sg13g2f_FILL8
XFILLER_42_1446 VDD VSS sg13g2f_FILL8
XFILLER_42_1454 VDD VSS sg13g2f_FILL8
XFILLER_42_1462 VDD VSS sg13g2f_FILL8
XFILLER_42_1470 VDD VSS sg13g2f_FILL8
XFILLER_42_1478 VDD VSS sg13g2f_FILL8
XFILLER_42_1486 VDD VSS sg13g2f_FILL8
XFILLER_42_1494 VDD VSS sg13g2f_FILL4
XFILLER_42_1505 VDD VSS sg13g2f_FILL8
XFILLER_42_1513 VDD VSS sg13g2f_FILL4
XFILLER_42_1531 VDD VSS sg13g2f_FILL8
XFILLER_42_1539 VDD VSS sg13g2f_FILL8
XFILLER_42_1547 VDD VSS sg13g2f_FILL4
XFILLER_43_1390 VDD VSS sg13g2f_FILL8
XFILLER_43_1398 VDD VSS sg13g2f_FILL8
XFILLER_43_1406 VDD VSS sg13g2f_FILL8
XFILLER_43_1414 VDD VSS sg13g2f_FILL8
XFILLER_43_1422 VDD VSS sg13g2f_FILL8
XFILLER_43_1430 VDD VSS sg13g2f_FILL8
XFILLER_43_1438 VDD VSS sg13g2f_FILL8
XFILLER_43_1446 VDD VSS sg13g2f_FILL8
XFILLER_43_1454 VDD VSS sg13g2f_FILL8
XFILLER_43_1462 VDD VSS sg13g2f_FILL8
XFILLER_43_1470 VDD VSS sg13g2f_FILL8
XFILLER_43_1478 VDD VSS sg13g2f_FILL8
XFILLER_43_1486 VDD VSS sg13g2f_FILL8
XFILLER_43_1494 VDD VSS sg13g2f_FILL8
XFILLER_43_1502 VDD VSS sg13g2f_FILL8
XFILLER_43_1510 VDD VSS sg13g2f_FILL8
XFILLER_43_1529 VDD VSS sg13g2f_FILL8
XFILLER_43_1537 VDD VSS sg13g2f_FILL8
XFILLER_43_1545 VDD VSS sg13g2f_FILL4
XFILLER_43_1549 VDD VSS sg13g2f_FILL2
XFILLER_44_1390 VDD VSS sg13g2f_FILL8
XFILLER_44_1398 VDD VSS sg13g2f_FILL8
XFILLER_44_1406 VDD VSS sg13g2f_FILL8
XFILLER_44_1414 VDD VSS sg13g2f_FILL8
XFILLER_44_1422 VDD VSS sg13g2f_FILL8
XFILLER_44_1430 VDD VSS sg13g2f_FILL8
XFILLER_44_1438 VDD VSS sg13g2f_FILL8
XFILLER_44_1446 VDD VSS sg13g2f_FILL8
XFILLER_44_1454 VDD VSS sg13g2f_FILL8
XFILLER_44_1462 VDD VSS sg13g2f_FILL8
XFILLER_44_1470 VDD VSS sg13g2f_FILL8
XFILLER_44_1478 VDD VSS sg13g2f_FILL8
XFILLER_44_1486 VDD VSS sg13g2f_FILL8
XFILLER_44_1494 VDD VSS sg13g2f_FILL4
XFILLER_44_1547 VDD VSS sg13g2f_FILL4
XFILLER_45_1390 VDD VSS sg13g2f_FILL8
XFILLER_45_1398 VDD VSS sg13g2f_FILL8
XFILLER_45_1406 VDD VSS sg13g2f_FILL8
XFILLER_45_1414 VDD VSS sg13g2f_FILL8
XFILLER_45_1422 VDD VSS sg13g2f_FILL8
XFILLER_45_1430 VDD VSS sg13g2f_FILL8
XFILLER_45_1438 VDD VSS sg13g2f_FILL8
XFILLER_45_1446 VDD VSS sg13g2f_FILL8
XFILLER_45_1454 VDD VSS sg13g2f_FILL8
XFILLER_45_1462 VDD VSS sg13g2f_FILL8
XFILLER_45_1470 VDD VSS sg13g2f_FILL8
XFILLER_45_1478 VDD VSS sg13g2f_FILL8
XFILLER_45_1486 VDD VSS sg13g2f_FILL8
XFILLER_45_1494 VDD VSS sg13g2f_FILL8
XFILLER_45_1502 VDD VSS sg13g2f_FILL8
XFILLER_45_1510 VDD VSS sg13g2f_FILL8
XFILLER_45_1529 VDD VSS sg13g2f_FILL8
XFILLER_45_1537 VDD VSS sg13g2f_FILL8
XFILLER_45_1545 VDD VSS sg13g2f_FILL4
XFILLER_45_1549 VDD VSS sg13g2f_FILL2
XFILLER_46_1390 VDD VSS sg13g2f_FILL8
XFILLER_46_1398 VDD VSS sg13g2f_FILL8
XFILLER_46_1406 VDD VSS sg13g2f_FILL8
XFILLER_46_1414 VDD VSS sg13g2f_FILL8
XFILLER_46_1422 VDD VSS sg13g2f_FILL8
XFILLER_46_1430 VDD VSS sg13g2f_FILL8
XFILLER_46_1438 VDD VSS sg13g2f_FILL8
XFILLER_46_1446 VDD VSS sg13g2f_FILL8
XFILLER_46_1454 VDD VSS sg13g2f_FILL8
XFILLER_46_1462 VDD VSS sg13g2f_FILL8
XFILLER_46_1470 VDD VSS sg13g2f_FILL8
XFILLER_46_1478 VDD VSS sg13g2f_FILL8
XFILLER_46_1486 VDD VSS sg13g2f_FILL8
XFILLER_46_1494 VDD VSS sg13g2f_FILL4
XFILLER_46_1505 VDD VSS sg13g2f_FILL8
XFILLER_46_1513 VDD VSS sg13g2f_FILL4
XFILLER_46_1517 VDD VSS sg13g2f_FILL1
XFILLER_46_1537 VDD VSS sg13g2f_FILL8
XFILLER_46_1545 VDD VSS sg13g2f_FILL4
XFILLER_46_1549 VDD VSS sg13g2f_FILL2
XFILLER_47_1390 VDD VSS sg13g2f_FILL8
XFILLER_47_1398 VDD VSS sg13g2f_FILL8
XFILLER_47_1406 VDD VSS sg13g2f_FILL8
XFILLER_47_1414 VDD VSS sg13g2f_FILL8
XFILLER_47_1422 VDD VSS sg13g2f_FILL8
XFILLER_47_1430 VDD VSS sg13g2f_FILL8
XFILLER_47_1438 VDD VSS sg13g2f_FILL8
XFILLER_47_1446 VDD VSS sg13g2f_FILL8
XFILLER_47_1454 VDD VSS sg13g2f_FILL8
XFILLER_47_1462 VDD VSS sg13g2f_FILL8
XFILLER_47_1470 VDD VSS sg13g2f_FILL8
XFILLER_47_1478 VDD VSS sg13g2f_FILL8
XFILLER_47_1486 VDD VSS sg13g2f_FILL8
XFILLER_47_1494 VDD VSS sg13g2f_FILL8
XFILLER_47_1502 VDD VSS sg13g2f_FILL4
XFILLER_47_1506 VDD VSS sg13g2f_FILL1
XFILLER_47_1534 VDD VSS sg13g2f_FILL8
XFILLER_47_1542 VDD VSS sg13g2f_FILL8
XFILLER_47_1550 VDD VSS sg13g2f_FILL1
XFILLER_48_1390 VDD VSS sg13g2f_FILL8
XFILLER_48_1398 VDD VSS sg13g2f_FILL8
XFILLER_48_1406 VDD VSS sg13g2f_FILL8
XFILLER_48_1414 VDD VSS sg13g2f_FILL8
XFILLER_48_1422 VDD VSS sg13g2f_FILL8
XFILLER_48_1430 VDD VSS sg13g2f_FILL8
XFILLER_48_1438 VDD VSS sg13g2f_FILL8
XFILLER_48_1446 VDD VSS sg13g2f_FILL8
XFILLER_48_1454 VDD VSS sg13g2f_FILL8
XFILLER_48_1462 VDD VSS sg13g2f_FILL8
XFILLER_48_1470 VDD VSS sg13g2f_FILL8
XFILLER_48_1478 VDD VSS sg13g2f_FILL8
XFILLER_48_1486 VDD VSS sg13g2f_FILL8
XFILLER_48_1494 VDD VSS sg13g2f_FILL4
XFILLER_48_1505 VDD VSS sg13g2f_FILL8
XFILLER_48_1513 VDD VSS sg13g2f_FILL4
XFILLER_48_1517 VDD VSS sg13g2f_FILL1
XFILLER_48_1529 VDD VSS sg13g2f_FILL8
XFILLER_48_1537 VDD VSS sg13g2f_FILL8
XFILLER_48_1545 VDD VSS sg13g2f_FILL4
XFILLER_48_1549 VDD VSS sg13g2f_FILL2
XFILLER_49_1390 VDD VSS sg13g2f_FILL8
XFILLER_49_1398 VDD VSS sg13g2f_FILL8
XFILLER_49_1406 VDD VSS sg13g2f_FILL8
XFILLER_49_1414 VDD VSS sg13g2f_FILL8
XFILLER_49_1422 VDD VSS sg13g2f_FILL8
XFILLER_49_1430 VDD VSS sg13g2f_FILL8
XFILLER_49_1438 VDD VSS sg13g2f_FILL8
XFILLER_49_1446 VDD VSS sg13g2f_FILL8
XFILLER_49_1454 VDD VSS sg13g2f_FILL8
XFILLER_49_1462 VDD VSS sg13g2f_FILL8
XFILLER_49_1470 VDD VSS sg13g2f_FILL8
XFILLER_49_1478 VDD VSS sg13g2f_FILL8
XFILLER_49_1486 VDD VSS sg13g2f_FILL8
XFILLER_49_1494 VDD VSS sg13g2f_FILL8
XFILLER_49_1502 VDD VSS sg13g2f_FILL8
XFILLER_49_1510 VDD VSS sg13g2f_FILL8
XFILLER_49_1518 VDD VSS sg13g2f_FILL8
XFILLER_49_1526 VDD VSS sg13g2f_FILL8
XFILLER_49_1534 VDD VSS sg13g2f_FILL8
XFILLER_49_1542 VDD VSS sg13g2f_FILL8
XFILLER_49_1550 VDD VSS sg13g2f_FILL1
XFILLER_50_1390 VDD VSS sg13g2f_FILL8
XFILLER_50_1398 VDD VSS sg13g2f_FILL8
XFILLER_50_1406 VDD VSS sg13g2f_FILL8
XFILLER_50_1414 VDD VSS sg13g2f_FILL8
XFILLER_50_1422 VDD VSS sg13g2f_FILL8
XFILLER_50_1430 VDD VSS sg13g2f_FILL8
XFILLER_50_1438 VDD VSS sg13g2f_FILL8
XFILLER_50_1446 VDD VSS sg13g2f_FILL8
XFILLER_50_1454 VDD VSS sg13g2f_FILL8
XFILLER_50_1462 VDD VSS sg13g2f_FILL8
XFILLER_50_1470 VDD VSS sg13g2f_FILL8
XFILLER_50_1478 VDD VSS sg13g2f_FILL8
XFILLER_50_1486 VDD VSS sg13g2f_FILL8
XFILLER_50_1494 VDD VSS sg13g2f_FILL4
XFILLER_50_1505 VDD VSS sg13g2f_FILL8
XFILLER_50_1513 VDD VSS sg13g2f_FILL8
XFILLER_50_1521 VDD VSS sg13g2f_FILL8
XFILLER_50_1529 VDD VSS sg13g2f_FILL8
XFILLER_50_1537 VDD VSS sg13g2f_FILL8
XFILLER_50_1545 VDD VSS sg13g2f_FILL4
XFILLER_50_1549 VDD VSS sg13g2f_FILL2
XFILLER_51_1390 VDD VSS sg13g2f_FILL8
XFILLER_51_1398 VDD VSS sg13g2f_FILL8
XFILLER_51_1406 VDD VSS sg13g2f_FILL8
XFILLER_51_1414 VDD VSS sg13g2f_FILL8
XFILLER_51_1422 VDD VSS sg13g2f_FILL8
XFILLER_51_1430 VDD VSS sg13g2f_FILL8
XFILLER_51_1438 VDD VSS sg13g2f_FILL8
XFILLER_51_1446 VDD VSS sg13g2f_FILL8
XFILLER_51_1454 VDD VSS sg13g2f_FILL8
XFILLER_51_1462 VDD VSS sg13g2f_FILL8
XFILLER_51_1470 VDD VSS sg13g2f_FILL8
XFILLER_51_1478 VDD VSS sg13g2f_FILL8
XFILLER_51_1486 VDD VSS sg13g2f_FILL8
XFILLER_51_1494 VDD VSS sg13g2f_FILL8
XFILLER_51_1502 VDD VSS sg13g2f_FILL8
XFILLER_51_1533 VDD VSS sg13g2f_FILL8
XFILLER_51_1541 VDD VSS sg13g2f_FILL8
XFILLER_51_1549 VDD VSS sg13g2f_FILL2
XFILLER_52_1390 VDD VSS sg13g2f_FILL8
XFILLER_52_1398 VDD VSS sg13g2f_FILL8
XFILLER_52_1406 VDD VSS sg13g2f_FILL8
XFILLER_52_1414 VDD VSS sg13g2f_FILL8
XFILLER_52_1422 VDD VSS sg13g2f_FILL8
XFILLER_52_1430 VDD VSS sg13g2f_FILL8
XFILLER_52_1438 VDD VSS sg13g2f_FILL8
XFILLER_52_1446 VDD VSS sg13g2f_FILL8
XFILLER_52_1454 VDD VSS sg13g2f_FILL8
XFILLER_52_1462 VDD VSS sg13g2f_FILL8
XFILLER_52_1470 VDD VSS sg13g2f_FILL8
XFILLER_52_1478 VDD VSS sg13g2f_FILL8
XFILLER_52_1486 VDD VSS sg13g2f_FILL8
XFILLER_52_1494 VDD VSS sg13g2f_FILL1
XFILLER_52_1502 VDD VSS sg13g2f_FILL8
XFILLER_52_1510 VDD VSS sg13g2f_FILL8
XFILLER_52_1518 VDD VSS sg13g2f_FILL8
XFILLER_52_1526 VDD VSS sg13g2f_FILL8
XFILLER_52_1534 VDD VSS sg13g2f_FILL8
XFILLER_52_1542 VDD VSS sg13g2f_FILL8
XFILLER_52_1550 VDD VSS sg13g2f_FILL1
.ENDS SARADC
* CDL Netlist generated by OpenROAD

*.BUSDELIMITER [

.SUBCKT SPI CEB CLK DATA DOUT_DAT DOUT_EN RD[0] RD[10] RD[11]
+ RD[12] RD[13] RD[14] RD[15] RD[16] RD[17] RD[18] RD[19] RD[1]
+ RD[20] RD[21] RD[22] RD[23] RD[24] RD[25] RD[26] RD[27] RD[28]
+ RD[29] RD[2] RD[30] RD[31] RD[32] RD[33] RD[34] RD[35] RD[36]
+ RD[37] RD[38] RD[39] RD[3] RD[40] RD[41] RD[42] RD[43] RD[44]
+ RD[45] RD[46] RD[47] RD[4] RD[5] RD[6] RD[7] RD[8] RD[9] RST
+ R[0] R[10] R[11] R[12] R[13] R[14] R[15] R[16] R[17] R[18]
+ R[19] R[1] R[20] R[21] R[22] R[23] R[24] R[25] R[26] R[27]
+ R[28] R[29] R[2] R[30] R[31] R[32] R[33] R[34] R[35] R[36]
+ R[37] R[38] R[39] R[3] R[40] R[41] R[42] R[43] R[44] R[45]
+ R[46] R[47] R[48] R[49] R[4] R[50] R[51] R[52] R[53] R[54]
+ R[55] R[56] R[57] R[58] R[59] R[5] R[60] R[61] R[62] R[63]
+ R[6] R[7] R[8] R[9] VSS VDD
Xins_223_ R[42] raddr\[2\] ins_124_ VDD VSS ins_036_ sg13g2_MUX2D1
Xins_224_ R[43] sft_reg\[3\] ins_124_ VDD VSS ins_037_ sg13g2_MUX2D1
Xins_225_ R[44] sft_reg\[4\] ins_124_ VDD VSS ins_038_ sg13g2_MUX2D1
Xins_226_ R[45] sft_reg\[5\] ins_124_ VDD VSS ins_039_ sg13g2_MUX2D1
Xins_227_ R[46] sft_reg\[6\] ins_124_ VDD VSS ins_040_ sg13g2_MUX2D1
Xins_228_ R[47] sft_reg\[7\] ins_124_ VDD VSS ins_041_ sg13g2_MUX2D1
Xins_229_ addr\[0\] addr\[1\] VDD VSS ins_125_ sg13g2_NR2D1
Xins_230_ ins_110_ ins_125_ VDD VSS ins_126_ sg13g2_AN2D1
Xins_231_ ins_121_ ins_126_ VDD VSS ins_127_ sg13g2_AN2D1
Xins_232_ R[0] raddr\[0\] ins_127_ VDD VSS ins_042_ sg13g2_MUX2D1
Xins_233_ R[1] raddr\[1\] ins_127_ VDD VSS ins_043_ sg13g2_MUX2D1
Xins_234_ R[2] raddr\[2\] ins_127_ VDD VSS ins_044_ sg13g2_MUX2D1
Xins_235_ R[3] sft_reg\[3\] ins_127_ VDD VSS ins_045_ sg13g2_MUX2D1
Xins_236_ R[4] sft_reg\[4\] ins_127_ VDD VSS ins_046_ sg13g2_MUX2D1
Xins_237_ R[5] sft_reg\[5\] ins_127_ VDD VSS ins_047_ sg13g2_MUX2D1
Xins_238_ R[6] sft_reg\[6\] ins_127_ VDD VSS ins_048_ sg13g2_MUX2D1
Xins_239_ R[7] sft_reg\[7\] ins_127_ VDD VSS ins_049_ sg13g2_MUX2D1
Xins_240_ ins_108_ addr\[1\] ins_110_ VDD VSS ins_128_ sg13g2_ND3D1
Xins_241_ ins_122_ ins_128_ VDD VSS ins_129_ sg13g2_NR2D1
Xins_242_ R[16] raddr\[0\] ins_129_ VDD VSS ins_050_ sg13g2_MUX2D1
Xins_243_ R[17] raddr\[1\] ins_129_ VDD VSS ins_051_ sg13g2_MUX2D1
Xins_244_ R[18] raddr\[2\] ins_129_ VDD VSS ins_052_ sg13g2_MUX2D1
Xins_245_ R[19] sft_reg\[3\] ins_129_ VDD VSS ins_053_ sg13g2_MUX2D1
Xins_246_ R[20] sft_reg\[4\] ins_129_ VDD VSS ins_054_ sg13g2_MUX2D1
Xins_247_ R[21] sft_reg\[5\] ins_129_ VDD VSS ins_055_ sg13g2_MUX2D1
Xins_248_ R[22] sft_reg\[6\] ins_129_ VDD VSS ins_056_ sg13g2_MUX2D1
Xins_249_ R[23] sft_reg\[7\] ins_129_ VDD VSS ins_057_ sg13g2_MUX2D1
Xins_250_ addr\[0\] addr\[1\] VDD VSS ins_130_ sg13g2_AN2D1
Xins_251_ addr\[2\] ins_121_ ins_130_ VDD VSS ins_131_ sg13g2_ND3D1
Xins_252_ raddr\[0\] R[56] ins_131_ VDD VSS ins_058_ sg13g2_MUX2D1
Xins_253_ raddr\[1\] R[57] ins_131_ VDD VSS ins_059_ sg13g2_MUX2D1
Xins_254_ raddr\[2\] R[58] ins_131_ VDD VSS ins_060_ sg13g2_MUX2D1
Xins_255_ sft_reg\[3\] R[59] ins_131_ VDD VSS ins_061_ sg13g2_MUX2D1
Xins_256_ sft_reg\[4\] R[60] ins_131_ VDD VSS ins_062_ sg13g2_MUX2D1
Xins_257_ sft_reg\[5\] R[61] ins_131_ VDD VSS ins_063_ sg13g2_MUX2D1
Xins_258_ sft_reg\[6\] R[62] ins_131_ VDD VSS ins_064_ sg13g2_MUX2D1
Xins_259_ sft_reg\[7\] R[63] ins_131_ VDD VSS ins_065_ sg13g2_MUX2D1
Xins_260_ genblk1.counter\[18\] genblk1.counter\[19\] VDD
+ VSS ins_132_ sg13g2_NR2D1
Xins_261_ genblk1.counter\[17\] genblk1.counter\[20\] VDD
+ VSS ins_133_ sg13g2_NR2D1
Xins_262_ genblk1.counter\[14\] genblk1.counter\[15\] VDD
+ VSS ins_134_ sg13g2_NR2D1
Xins_263_ genblk1.counter\[13\] genblk1.counter\[16\] VDD
+ VSS ins_135_ sg13g2_NR2D1
Xins_264_ ins_132_ ins_133_ ins_134_ ins_135_ VDD VSS ins_136_
+ sg13g2_ND4D1
Xins_265_ re ins_136_ VDD VSS ins_137_ sg13g2_ND2D1
Xins_266_ ins_137_ eno VSS VDD sg13g2_INVD1
Xins_267_ addr\[0\] ins_109_ ins_110_ VDD VSS ins_138_ sg13g2_ND3D1
Xins_268_ addr\[0\] ins_109_ ins_110_ RD[8] VDD VSS ins_139_
+ sg13g2_ND4D1
Xins_269_ ins_110_ RD[0] ins_125_ VDD VSS ins_140_ sg13g2_ND3D1
Xins_270_ addr\[2\] RD[32] ins_125_ VDD VSS ins_141_ sg13g2_ND3D1
Xins_271_ addr\[0\] ins_109_ addr\[2\] RD[40] VDD VSS ins_142_
+ sg13g2_ND4D1
Xins_272_ ins_108_ addr\[1\] ins_110_ RD[16] VDD VSS ins_143_
+ sg13g2_ND4D1
Xins_273_ ins_110_ ins_130_ VDD VSS ins_144_ sg13g2_AN2D1
Xins_274_ ins_110_ RD[24] ins_130_ VDD VSS ins_145_ sg13g2_ND3D1
Xins_275_ ins_139_ ins_140_ ins_143_ ins_145_ VDD VSS ins_146_
+ sg13g2_ND4D1
Xins_276_ encap ins_141_ ins_142_ VDD VSS ins_147_ sg13g2_ND3D1
Xins_277_ bus_cap\[0\] ins_137_ encap VDD VSS ins_148_ sg13g2_AO21D1
Xins_278_ ins_146_ ins_147_ ins_148_ VDD VSS ins_066_ sg13g2_OA21D1
Xins_279_ bus_cap\[0\] bus_cap\[1\] ins_137_ VDD VSS ins_149_
+ sg13g2_MUX2D1
Xins_280_ ins_108_ addr\[1\] ins_110_ RD[17] VDD VSS ins_150_
+ sg13g2_ND4D1
Xins_281_ ins_110_ RD[1] ins_125_ VDD VSS ins_151_ sg13g2_ND3D1
Xins_282_ ins_150_ ins_151_ VDD VSS ins_152_ sg13g2_AN2D1
Xins_283_ addr\[2\] RD[33] ins_125_ VDD VSS ins_153_ sg13g2_ND3D1
Xins_284_ addr\[0\] ins_109_ ins_110_ RD[9] VDD VSS ins_154_
+ sg13g2_ND4D1
Xins_285_ ins_153_ ins_154_ VDD VSS ins_155_ sg13g2_AN2D1
Xins_286_ addr\[0\] ins_109_ addr\[2\] RD[41] VDD VSS ins_156_
+ sg13g2_ND4D1
Xins_287_ ins_110_ RD[25] ins_130_ VDD VSS ins_157_ sg13g2_ND3D1
Xins_288_ ins_152_ ins_155_ ins_156_ ins_157_ VDD VSS ins_158_
+ sg13g2_ND4D1
Xins_289_ ins_149_ ins_158_ encap VDD VSS ins_067_ sg13g2_MUX2D1
Xins_290_ bus_cap\[1\] bus_cap\[2\] ins_137_ VDD VSS ins_159_
+ sg13g2_MUX2D1
Xins_291_ addr\[2\] RD[34] ins_125_ VDD VSS ins_160_ sg13g2_ND3D1
Xins_292_ addr\[0\] ins_109_ ins_110_ RD[10] VDD VSS ins_161_
+ sg13g2_ND4D1
Xins_293_ ins_160_ ins_161_ VDD VSS ins_162_ sg13g2_ND2D1
Xins_294_ ins_110_ RD[26] ins_130_ VDD VSS ins_163_ sg13g2_ND3D1
Xins_295_ ins_108_ addr\[1\] ins_110_ RD[18] VDD VSS ins_164_
+ sg13g2_ND4D1
Xins_296_ ins_110_ RD[2] ins_125_ VDD VSS ins_165_ sg13g2_ND3D1
Xins_297_ addr\[0\] ins_109_ addr\[2\] RD[42] VDD VSS ins_166_
+ sg13g2_ND4D1
Xins_298_ ins_163_ ins_164_ ins_165_ ins_166_ VDD VSS ins_167_
+ sg13g2_ND4D1
Xins_299_ ins_162_ ins_167_ VDD VSS ins_168_ sg13g2_OR2D1
Xins_300_ ins_159_ ins_168_ encap VDD VSS ins_068_ sg13g2_MUX2D1
Xins_301_ bus_cap\[2\] bus_cap\[3\] ins_137_ VDD VSS ins_169_
+ sg13g2_MUX2D1
Xins_302_ addr\[0\] ins_109_ ins_110_ RD[11] VDD VSS ins_170_
+ sg13g2_ND4D1
Xins_303_ ins_110_ RD[27] ins_130_ VDD VSS ins_171_ sg13g2_ND3D1
Xins_304_ ins_170_ ins_171_ VDD VSS ins_172_ sg13g2_ND2D1
Xins_305_ ins_110_ RD[3] ins_125_ VDD VSS ins_173_ sg13g2_ND3D1
Xins_306_ ins_108_ addr\[1\] ins_110_ RD[19] VDD VSS ins_174_
+ sg13g2_ND4D1
Xins_307_ addr\[2\] RD[35] ins_125_ VDD VSS ins_175_ sg13g2_ND3D1
Xins_308_ addr\[0\] ins_109_ addr\[2\] RD[43] VDD VSS ins_176_
+ sg13g2_ND4D1
Xins_309_ ins_173_ ins_174_ ins_175_ ins_176_ VDD VSS ins_177_
+ sg13g2_ND4D1
Xins_310_ ins_172_ ins_177_ VDD VSS ins_178_ sg13g2_OR2D1
Xins_311_ ins_169_ ins_178_ encap VDD VSS ins_069_ sg13g2_MUX2D1
Xins_312_ bus_cap\[3\] bus_cap\[4\] ins_137_ VDD VSS ins_179_
+ sg13g2_MUX2D1
Xins_313_ addr\[0\] ins_109_ ins_110_ RD[12] VDD VSS ins_180_
+ sg13g2_ND4D1
Xins_314_ ins_108_ addr\[1\] ins_110_ RD[20] VDD VSS ins_181_
+ sg13g2_ND4D1
Xins_315_ ins_180_ ins_181_ VDD VSS ins_182_ sg13g2_ND2D1
Xins_316_ ins_110_ RD[4] ins_125_ VDD VSS ins_183_ sg13g2_ND3D1
Xins_317_ ins_110_ RD[28] ins_130_ VDD VSS ins_184_ sg13g2_ND3D1
Xins_318_ addr\[2\] RD[36] ins_125_ VDD VSS ins_185_ sg13g2_ND3D1
Xins_319_ addr\[0\] ins_109_ addr\[2\] RD[44] VDD VSS ins_186_
+ sg13g2_ND4D1
Xins_320_ ins_183_ ins_184_ ins_185_ ins_186_ VDD VSS ins_187_
+ sg13g2_ND4D1
Xins_321_ ins_182_ ins_187_ VDD VSS ins_188_ sg13g2_OR2D1
Xins_322_ ins_179_ ins_188_ encap VDD VSS ins_070_ sg13g2_MUX2D1
Xins_323_ bus_cap\[4\] bus_cap\[5\] ins_137_ VDD VSS ins_189_
+ sg13g2_MUX2D1
Xins_324_ addr\[0\] ins_109_ ins_110_ RD[13] VDD VSS ins_190_
+ sg13g2_ND4D1
Xins_325_ ins_110_ RD[29] ins_130_ VDD VSS ins_191_ sg13g2_ND3D1
Xins_326_ ins_190_ ins_191_ VDD VSS ins_192_ sg13g2_ND2D1
Xins_327_ ins_110_ RD[5] ins_125_ VDD VSS ins_193_ sg13g2_ND3D1
Xins_328_ ins_108_ addr\[1\] ins_110_ RD[21] VDD VSS ins_194_
+ sg13g2_ND4D1
Xins_329_ addr\[2\] RD[37] ins_125_ VDD VSS ins_195_ sg13g2_ND3D1
Xins_330_ addr\[0\] ins_109_ addr\[2\] RD[45] VDD VSS ins_196_
+ sg13g2_ND4D1
Xins_331_ ins_193_ ins_194_ ins_195_ ins_196_ VDD VSS ins_197_
+ sg13g2_ND4D1
Xins_332_ ins_192_ ins_197_ VDD VSS ins_198_ sg13g2_OR2D1
Xins_333_ ins_189_ ins_198_ encap VDD VSS ins_071_ sg13g2_MUX2D1
Xins_334_ bus_cap\[5\] bus_cap\[6\] ins_137_ VDD VSS ins_199_
+ sg13g2_MUX2D1
Xins_335_ ins_110_ RD[6] ins_125_ VDD VSS ins_200_ sg13g2_ND3D1
Xins_336_ ins_108_ addr\[1\] ins_110_ RD[22] VDD VSS ins_201_
+ sg13g2_ND4D1
Xins_337_ ins_200_ ins_201_ VDD VSS ins_202_ sg13g2_AN2D1
Xins_338_ addr\[0\] ins_109_ addr\[2\] RD[46] VDD VSS ins_203_
+ sg13g2_ND4D1
Xins_339_ ins_110_ RD[30] ins_130_ VDD VSS ins_204_ sg13g2_ND3D1
Xins_340_ addr\[2\] RD[38] ins_125_ VDD VSS ins_205_ sg13g2_ND3D1
Xins_341_ addr\[0\] ins_109_ ins_110_ RD[14] VDD VSS ins_206_
+ sg13g2_ND4D1
Xins_342_ ins_205_ ins_206_ VDD VSS ins_207_ sg13g2_AN2D1
Xins_343_ ins_202_ ins_203_ ins_204_ ins_207_ VDD VSS ins_208_
+ sg13g2_ND4D1
Xins_344_ ins_199_ ins_208_ encap VDD VSS ins_072_ sg13g2_MUX2D1
Xins_345_ bus_cap\[6\] bus_cap\[7\] ins_137_ VDD VSS ins_209_
+ sg13g2_MUX2D1
Xins_346_ addr\[2\] RD[39] ins_125_ VDD VSS ins_210_ sg13g2_ND3D1
Xins_347_ addr\[0\] ins_109_ ins_110_ RD[15] VDD VSS ins_211_
+ sg13g2_ND4D1
Xins_348_ ins_108_ addr\[1\] ins_110_ RD[23] VDD VSS ins_212_
+ sg13g2_ND4D1
Xins_349_ ins_110_ RD[7] ins_125_ VDD VSS ins_213_ sg13g2_ND3D1
Xins_350_ ins_212_ ins_213_ VDD VSS ins_214_ sg13g2_AN2D1
Xins_351_ ins_110_ RD[31] ins_130_ VDD VSS ins_215_ sg13g2_ND3D1
Xins_352_ addr\[0\] ins_109_ addr\[2\] RD[47] VDD VSS ins_216_
+ sg13g2_ND4D1
Xins_353_ ins_211_ ins_216_ VDD VSS ins_217_ sg13g2_AN2D1
Xins_354_ ins_210_ ins_214_ ins_215_ ins_217_ VDD VSS ins_218_
+ sg13g2_ND4D1
Xins_355_ ins_209_ ins_218_ encap VDD VSS ins_073_ sg13g2_MUX2D1
Xins_356_ ins_108_ addr\[1\] addr\[2\] ins_121_ VDD VSS ins_219_
+ sg13g2_ND4D1
Xins_357_ raddr\[0\] R[48] ins_219_ VDD VSS ins_074_ sg13g2_MUX2D1
Xins_358_ raddr\[1\] R[49] ins_219_ VDD VSS ins_075_ sg13g2_MUX2D1
Xins_359_ raddr\[2\] R[50] ins_219_ VDD VSS ins_076_ sg13g2_MUX2D1
Xins_360_ sft_reg\[3\] R[51] ins_219_ VDD VSS ins_077_ sg13g2_MUX2D1
Xins_361_ sft_reg\[4\] R[52] ins_219_ VDD VSS ins_078_ sg13g2_MUX2D1
Xins_362_ sft_reg\[5\] R[53] ins_219_ VDD VSS ins_079_ sg13g2_MUX2D1
Xins_363_ sft_reg\[6\] R[54] ins_219_ VDD VSS ins_080_ sg13g2_MUX2D1
Xins_364_ sft_reg\[7\] R[55] ins_219_ VDD VSS ins_081_ sg13g2_MUX2D1
Xins_365_ CEB ins_021_ VDD VSS ins_011_ sg13g2_NR2D1
Xins_366_ we DATA ins_011_ VDD VSS ins_082_ sg13g2_MUX2D1
Xins_367_ addr\[2\] ins_121_ ins_125_ VDD VSS ins_220_ sg13g2_ND3D1
Xins_368_ raddr\[0\] R[32] ins_220_ VDD VSS ins_083_ sg13g2_MUX2D1
Xins_369_ raddr\[1\] R[33] ins_220_ VDD VSS ins_084_ sg13g2_MUX2D1
Xins_370_ raddr\[2\] R[34] ins_220_ VDD VSS ins_085_ sg13g2_MUX2D1
Xins_371_ sft_reg\[3\] R[35] ins_220_ VDD VSS ins_086_ sg13g2_MUX2D1
Xins_372_ sft_reg\[4\] R[36] ins_220_ VDD VSS ins_087_ sg13g2_MUX2D1
Xins_373_ sft_reg\[5\] R[37] ins_220_ VDD VSS ins_088_ sg13g2_MUX2D1
Xins_374_ sft_reg\[6\] R[38] ins_220_ VDD VSS ins_089_ sg13g2_MUX2D1
Xins_375_ sft_reg\[7\] R[39] ins_220_ VDD VSS ins_090_ sg13g2_MUX2D1
Xins_376_ ins_121_ ins_144_ VDD VSS ins_221_ sg13g2_AN2D1
Xins_377_ R[24] raddr\[0\] ins_221_ VDD VSS ins_091_ sg13g2_MUX2D1
Xins_378_ R[25] raddr\[1\] ins_221_ VDD VSS ins_092_ sg13g2_MUX2D1
Xins_379_ R[26] raddr\[2\] ins_221_ VDD VSS ins_093_ sg13g2_MUX2D1
Xins_380_ R[27] sft_reg\[3\] ins_221_ VDD VSS ins_094_ sg13g2_MUX2D1
Xins_381_ R[28] sft_reg\[4\] ins_221_ VDD VSS ins_095_ sg13g2_MUX2D1
Xins_382_ R[29] sft_reg\[5\] ins_221_ VDD VSS ins_096_ sg13g2_MUX2D1
Xins_383_ R[30] sft_reg\[6\] ins_221_ VDD VSS ins_097_ sg13g2_MUX2D1
Xins_384_ R[31] sft_reg\[7\] ins_221_ VDD VSS ins_098_ sg13g2_MUX2D1
Xins_385_ ins_122_ ins_138_ VDD VSS ins_222_ sg13g2_NR2D1
Xins_386_ R[8] raddr\[0\] ins_222_ VDD VSS ins_099_ sg13g2_MUX2D1
Xins_387_ R[9] raddr\[1\] ins_222_ VDD VSS ins_100_ sg13g2_MUX2D1
Xins_388_ R[10] raddr\[2\] ins_222_ VDD VSS ins_101_ sg13g2_MUX2D1
Xins_389_ R[11] sft_reg\[3\] ins_222_ VDD VSS ins_102_ sg13g2_MUX2D1
Xins_390_ R[12] sft_reg\[4\] ins_222_ VDD VSS ins_103_ sg13g2_MUX2D1
Xins_391_ R[13] sft_reg\[5\] ins_222_ VDD VSS ins_104_ sg13g2_MUX2D1
Xins_392_ R[14] sft_reg\[6\] ins_222_ VDD VSS ins_105_ sg13g2_MUX2D1
Xins_393_ R[15] sft_reg\[7\] ins_222_ VDD VSS ins_106_ sg13g2_MUX2D1
Xins_394_ ins_022_ genblk1.counter\[1\] VDD VSS ins_013_ sg13g2_AN2D1
Xins_395_ re DATA ins_013_ VDD VSS ins_107_ sg13g2_MUX2D1
Xins_396_ ins_022_ genblk1.counter\[2\] VDD VSS ins_014_ sg13g2_AN2D1
Xins_397_ ins_022_ genblk1.counter\[3\] VDD VSS ins_015_ sg13g2_AN2D1
Xins_398_ ins_022_ genblk1.counter\[4\] VDD VSS ins_016_ sg13g2_AN2D1
Xins_399_ ins_022_ encap VDD VSS ins_017_ sg13g2_AN2D1
Xins_400_ ins_022_ genblk1.counter\[6\] VDD VSS ins_018_ sg13g2_AN2D1
Xins_401_ ins_022_ genblk1.counter\[7\] VDD VSS ins_019_ sg13g2_AN2D1
Xins_402_ ins_022_ genblk1.counter\[8\] VDD VSS ins_020_ sg13g2_AN2D1
Xins_403_ ins_022_ genblk1.counter\[9\] VDD VSS ins_001_ sg13g2_AN2D1
Xins_404_ ins_022_ genblk1.counter\[10\] VDD VSS ins_002_
+ sg13g2_AN2D1
Xins_405_ ins_022_ genblk1.counter\[11\] VDD VSS ins_003_
+ sg13g2_AN2D1
Xins_406_ ins_022_ genblk1.counter\[12\] VDD VSS ins_004_
+ sg13g2_AN2D1
Xins_407_ ins_022_ genblk1.counter\[13\] VDD VSS ins_005_
+ sg13g2_AN2D1
Xins_408_ ins_022_ genblk1.counter\[14\] VDD VSS ins_006_
+ sg13g2_AN2D1
Xins_409_ ins_022_ genblk1.counter\[15\] VDD VSS ins_007_
+ sg13g2_AN2D1
Xins_410_ ins_022_ genblk1.counter\[16\] VDD VSS ins_008_
+ sg13g2_AN2D1
Xins_411_ ins_022_ genblk1.counter\[17\] VDD VSS ins_009_
+ sg13g2_AN2D1
Xins_412_ ins_022_ genblk1.counter\[18\] VDD VSS ins_010_
+ sg13g2_AN2D1
Xins_413_ ins_022_ genblk1.counter\[19\] VDD VSS ins_012_
+ sg13g2_AN2D1
Xins_414_ bus_cap\[7\] eno VDD VSS ins_000_ sg13g2_AN2D1
Xins_415_ ins_022_ enoz VDD VSS DOUT_EN sg13g2_AN2D1
Xins_416_ CEB ins_022_ VSS VDD sg13g2_INVD1
Xins_417_ addr\[0\] ins_108_ VSS VDD sg13g2_INVD1
Xins_418_ addr\[1\] ins_109_ VSS VDD sg13g2_INVD1
Xins_419_ addr\[2\] ins_110_ VSS VDD sg13g2_INVD1
Xins_420_ genblk1.counter\[1\] ins_111_ VSS VDD sg13g2_INVD1
Xins_421_ genblk1.counter\[12\] ins_112_ VSS VDD sg13g2_INVD1
Xins_422_ genblk1.counter\[2\] genblk1.counter\[3\] VDD VSS
+ ins_113_ sg13g2_NR2D1
Xins_423_ genblk1.counter\[4\] encap VDD VSS ins_114_ sg13g2_NR2D1
Xins_424_ ins_021_ ins_111_ ins_113_ ins_114_ VDD VSS ins_115_
+ sg13g2_ND4D1
Xins_425_ genblk1.counter\[10\] genblk1.counter\[11\] VDD
+ VSS ins_116_ sg13g2_NR2D1
Xins_426_ genblk1.counter\[6\] genblk1.counter\[7\] VDD VSS
+ ins_117_ sg13g2_NR2D1
Xins_427_ genblk1.counter\[8\] genblk1.counter\[9\] VDD VSS
+ ins_118_ sg13g2_NR2D1
Xins_428_ ins_112_ ins_116_ ins_117_ ins_118_ VDD VSS ins_119_
+ sg13g2_ND4D1
Xins_429_ ins_115_ ins_119_ ins_022_ VDD VSS ins_120_ sg13g2_OAI21D1
Xins_430_ DATA raddr\[0\] ins_120_ VDD VSS ins_023_ sg13g2_MUX2D1
Xins_431_ raddr\[0\] raddr\[1\] ins_120_ VDD VSS ins_024_
+ sg13g2_MUX2D1
Xins_432_ raddr\[1\] raddr\[2\] ins_120_ VDD VSS ins_025_
+ sg13g2_MUX2D1
Xins_433_ raddr\[2\] sft_reg\[3\] ins_120_ VDD VSS ins_026_
+ sg13g2_MUX2D1
Xins_434_ sft_reg\[3\] sft_reg\[4\] ins_120_ VDD VSS ins_027_
+ sg13g2_MUX2D1
Xins_435_ sft_reg\[4\] sft_reg\[5\] ins_120_ VDD VSS ins_028_
+ sg13g2_MUX2D1
Xins_436_ sft_reg\[5\] sft_reg\[6\] ins_120_ VDD VSS ins_029_
+ sg13g2_MUX2D1
Xins_437_ sft_reg\[6\] sft_reg\[7\] ins_120_ VDD VSS ins_030_
+ sg13g2_MUX2D1
Xins_438_ sft_reg\[7\] addr\[0\] ins_120_ VDD VSS ins_031_
+ sg13g2_MUX2D1
Xins_439_ addr\[0\] addr\[1\] ins_120_ VDD VSS ins_032_ sg13g2_MUX2D1
Xins_440_ addr\[1\] addr\[2\] ins_120_ VDD VSS ins_033_ sg13g2_MUX2D1
Xins_441_ we genblk1.counter\[13\] VDD VSS ins_121_ sg13g2_AN2D1
Xins_442_ we genblk1.counter\[13\] VDD VSS ins_122_ sg13g2_ND2D1
Xins_443_ addr\[0\] ins_109_ addr\[2\] VDD VSS ins_123_ sg13g2_ND3D1
Xins_444_ ins_122_ ins_123_ VDD VSS ins_124_ sg13g2_NR2D1
Xins_445_ R[40] raddr\[0\] ins_124_ VDD VSS ins_034_ sg13g2_MUX2D1
Xins_446_ R[41] raddr\[1\] ins_124_ VDD VSS ins_035_ sg13g2_MUX2D1
Xins_447_ RST clknet_3_2__leaf_CLK ins_023_ raddr\[0\] VDD
+ VSS sg13g2_DFCNQD1
Xins_448_ RST clknet_3_2__leaf_CLK ins_024_ raddr\[1\] VDD
+ VSS sg13g2_DFCNQD1
Xins_449_ RST clknet_3_2__leaf_CLK ins_025_ raddr\[2\] VDD
+ VSS sg13g2_DFCNQD1
Xins_450_ RST clknet_3_2__leaf_CLK ins_026_ sft_reg\[3\] VDD
+ VSS sg13g2_DFCNQD1
Xins_451_ RST clknet_3_2__leaf_CLK ins_027_ sft_reg\[4\] VDD
+ VSS sg13g2_DFCNQD1
Xins_452_ RST clknet_3_2__leaf_CLK ins_028_ sft_reg\[5\] VDD
+ VSS sg13g2_DFCNQD1
Xins_453_ RST clknet_3_0__leaf_CLK ins_029_ sft_reg\[6\] VDD
+ VSS sg13g2_DFCNQD1
Xins_454_ RST clknet_3_2__leaf_CLK ins_030_ sft_reg\[7\] VDD
+ VSS sg13g2_DFCNQD1
Xins_455_ RST clknet_3_3__leaf_CLK ins_031_ addr\[0\] VDD
+ VSS sg13g2_DFCNQD1
Xins_456_ RST clknet_3_3__leaf_CLK ins_032_ addr\[1\] VDD
+ VSS sg13g2_DFCNQD1
Xins_457_ RST clknet_3_3__leaf_CLK ins_033_ addr\[2\] VDD
+ VSS sg13g2_DFCNQD1
Xins_458_ RST clknet_3_0__leaf_CLK ins_034_ R[40] VDD VSS
+ sg13g2_DFCNQD1
Xins_459_ RST clknet_3_4__leaf_CLK ins_035_ R[41] VDD VSS
+ sg13g2_DFCNQD1
Xins_460_ RST clknet_3_0__leaf_CLK ins_036_ R[42] VDD VSS
+ sg13g2_DFCNQD1
Xins_461_ RST clknet_3_7__leaf_CLK ins_037_ R[43] VDD VSS
+ sg13g2_DFCNQD1
Xins_462_ RST clknet_3_3__leaf_CLK ins_038_ R[44] VDD VSS
+ sg13g2_DFCNQD1
Xins_463_ RST clknet_3_0__leaf_CLK ins_039_ R[45] VDD VSS
+ sg13g2_DFCNQD1
Xins_464_ RST clknet_3_3__leaf_CLK ins_040_ R[46] VDD VSS
+ sg13g2_DFCNQD1
Xins_465_ RST clknet_3_5__leaf_CLK ins_041_ R[47] VDD VSS
+ sg13g2_DFCNQD1
Xins_466_ RST clknet_3_4__leaf_CLK ins_042_ R[0] VDD VSS sg13g2_DFCNQD1
Xins_467_ RST clknet_3_5__leaf_CLK ins_043_ R[1] VDD VSS sg13g2_DFCNQD1
Xins_468_ RST clknet_3_0__leaf_CLK ins_044_ R[2] VDD VSS sg13g2_DFCNQD1
Xins_469_ RST clknet_3_5__leaf_CLK ins_045_ R[3] VDD VSS sg13g2_DFCNQD1
Xins_470_ RST clknet_3_5__leaf_CLK ins_046_ R[4] VDD VSS sg13g2_DFCNQD1
Xins_471_ RST clknet_3_1__leaf_CLK ins_047_ R[5] VDD VSS sg13g2_DFCNQD1
Xins_472_ RST clknet_3_1__leaf_CLK ins_048_ R[6] VDD VSS sg13g2_DFCNQD1
Xins_473_ RST clknet_3_5__leaf_CLK ins_049_ R[7] VDD VSS sg13g2_DFCNQD1
Xins_474_ RST clknet_3_2__leaf_CLK ins_050_ R[16] VDD VSS
+ sg13g2_DFCNQD1
Xins_475_ RST clknet_3_2__leaf_CLK ins_051_ R[17] VDD VSS
+ sg13g2_DFCNQD1
Xins_476_ RST clknet_3_6__leaf_CLK ins_052_ R[18] VDD VSS
+ sg13g2_DFCNQD1
Xins_477_ RST clknet_3_7__leaf_CLK ins_053_ R[19] VDD VSS
+ sg13g2_DFCNQD1
Xins_478_ RST clknet_3_6__leaf_CLK ins_054_ R[20] VDD VSS
+ sg13g2_DFCNQD1
Xins_479_ RST clknet_3_6__leaf_CLK ins_055_ R[21] VDD VSS
+ sg13g2_DFCNQD1
Xins_480_ RST clknet_3_7__leaf_CLK ins_056_ R[22] VDD VSS
+ sg13g2_DFCNQD1
Xins_481_ RST clknet_3_3__leaf_CLK ins_057_ R[23] VDD VSS
+ sg13g2_DFCNQD1
Xins_482_ RST clknet_3_0__leaf_CLK ins_058_ R[56] VDD VSS
+ sg13g2_DFCNQD1
Xins_483_ RST clknet_3_0__leaf_CLK ins_059_ R[57] VDD VSS
+ sg13g2_DFCNQD1
Xins_484_ RST clknet_3_5__leaf_CLK ins_060_ R[58] VDD VSS
+ sg13g2_DFCNQD1
Xins_485_ RST clknet_3_5__leaf_CLK ins_061_ R[59] VDD VSS
+ sg13g2_DFCNQD1
Xins_486_ RST clknet_3_0__leaf_CLK ins_062_ R[60] VDD VSS
+ sg13g2_DFCNQD1
Xins_487_ RST clknet_3_4__leaf_CLK ins_063_ R[61] VDD VSS
+ sg13g2_DFCNQD1
Xins_488_ RST clknet_3_1__leaf_CLK ins_064_ R[62] VDD VSS
+ sg13g2_DFCNQD1
Xins_489_ RST clknet_3_5__leaf_CLK ins_065_ R[63] VDD VSS
+ sg13g2_DFCNQD1
Xins_490_ RST clknet_3_4__leaf_CLK ins_066_ bus_cap\[0\] VDD
+ VSS sg13g2_DFCNQD1
Xins_491_ RST clknet_3_5__leaf_CLK ins_067_ bus_cap\[1\] VDD
+ VSS sg13g2_DFCNQD1
Xins_492_ RST clknet_3_7__leaf_CLK ins_068_ bus_cap\[2\] VDD
+ VSS sg13g2_DFCNQD1
Xins_493_ RST clknet_3_7__leaf_CLK ins_069_ bus_cap\[3\] VDD
+ VSS sg13g2_DFCNQD1
Xins_494_ RST clknet_3_7__leaf_CLK ins_070_ bus_cap\[4\] VDD
+ VSS sg13g2_DFCNQD1
Xins_495_ RST clknet_3_3__leaf_CLK ins_071_ bus_cap\[5\] VDD
+ VSS sg13g2_DFCNQD1
Xins_496_ RST clknet_3_3__leaf_CLK ins_072_ bus_cap\[6\] VDD
+ VSS sg13g2_DFCNQD1
Xins_497_ RST clknet_3_3__leaf_CLK ins_073_ bus_cap\[7\] VDD
+ VSS sg13g2_DFCNQD1
Xins_498_ RST clknet_3_0__leaf_CLK ins_074_ R[48] VDD VSS
+ sg13g2_DFCNQD1
Xins_499_ RST clknet_3_5__leaf_CLK ins_075_ R[49] VDD VSS
+ sg13g2_DFCNQD1
Xins_500_ RST clknet_3_5__leaf_CLK ins_076_ R[50] VDD VSS
+ sg13g2_DFCNQD1
Xins_501_ RST clknet_3_0__leaf_CLK ins_077_ R[51] VDD VSS
+ sg13g2_DFCNQD1
Xins_502_ RST clknet_3_1__leaf_CLK ins_078_ R[52] VDD VSS
+ sg13g2_DFCNQD1
Xins_503_ RST clknet_3_0__leaf_CLK ins_079_ R[53] VDD VSS
+ sg13g2_DFCNQD1
Xins_504_ RST clknet_3_5__leaf_CLK ins_080_ R[54] VDD VSS
+ sg13g2_DFCNQD1
Xins_505_ RST clknet_3_0__leaf_CLK ins_081_ R[55] VDD VSS
+ sg13g2_DFCNQD1
Xins_506_ RST clknet_3_6__leaf_CLK ins_082_ we VDD VSS sg13g2_DFCNQD1
Xins_507_ RST clknet_3_7__leaf_CLK ins_022_ ins_021_ VDD VSS
+ sg13g2_DFCNQD1
Xins_508_ RST clknet_3_6__leaf_CLK ins_011_ genblk1.counter\[1\]
+ VDD VSS sg13g2_DFCNQD1
Xins_509_ RST clknet_3_6__leaf_CLK ins_013_ genblk1.counter\[2\]
+ VDD VSS sg13g2_DFCNQD1
Xins_510_ RST clknet_3_7__leaf_CLK ins_014_ genblk1.counter\[3\]
+ VDD VSS sg13g2_DFCNQD1
Xins_511_ RST clknet_3_7__leaf_CLK ins_015_ genblk1.counter\[4\]
+ VDD VSS sg13g2_DFCNQD1
Xins_512_ RST clknet_3_7__leaf_CLK ins_016_ encap VDD VSS
+ sg13g2_DFCNQD1
Xins_513_ RST clknet_3_2__leaf_CLK ins_017_ genblk1.counter\[6\]
+ VDD VSS sg13g2_DFCNQD1
Xins_514_ RST clknet_3_2__leaf_CLK ins_018_ genblk1.counter\[7\]
+ VDD VSS sg13g2_DFCNQD1
Xins_515_ RST clknet_3_2__leaf_CLK ins_019_ genblk1.counter\[8\]
+ VDD VSS sg13g2_DFCNQD1
Xins_516_ RST clknet_3_2__leaf_CLK ins_020_ genblk1.counter\[9\]
+ VDD VSS sg13g2_DFCNQD1
Xins_517_ RST clknet_3_2__leaf_CLK ins_001_ genblk1.counter\[10\]
+ VDD VSS sg13g2_DFCNQD1
Xins_518_ RST clknet_3_3__leaf_CLK ins_002_ genblk1.counter\[11\]
+ VDD VSS sg13g2_DFCNQD1
Xins_519_ RST clknet_3_6__leaf_CLK ins_003_ genblk1.counter\[12\]
+ VDD VSS sg13g2_DFCNQD1
Xins_520_ RST clknet_3_3__leaf_CLK ins_004_ genblk1.counter\[13\]
+ VDD VSS sg13g2_DFCNQD1
Xins_521_ RST clknet_3_6__leaf_CLK ins_005_ genblk1.counter\[14\]
+ VDD VSS sg13g2_DFCNQD1
Xins_522_ RST clknet_3_6__leaf_CLK ins_006_ genblk1.counter\[15\]
+ VDD VSS sg13g2_DFCNQD1
Xins_523_ RST clknet_3_6__leaf_CLK ins_007_ genblk1.counter\[16\]
+ VDD VSS sg13g2_DFCNQD1
Xins_524_ RST clknet_3_6__leaf_CLK ins_008_ genblk1.counter\[17\]
+ VDD VSS sg13g2_DFCNQD1
Xins_525_ RST clknet_3_7__leaf_CLK ins_009_ genblk1.counter\[18\]
+ VDD VSS sg13g2_DFCNQD1
Xins_526_ RST clknet_3_7__leaf_CLK ins_010_ genblk1.counter\[19\]
+ VDD VSS sg13g2_DFCNQD1
Xins_527_ RST clknet_3_7__leaf_CLK ins_012_ genblk1.counter\[20\]
+ VDD VSS sg13g2_DFCNQD1
Xins_528_ RST clknet_3_3__leaf_CLK eno enoz VDD VSS sg13g2_DFCNQD1
Xins_529_ RST clknet_3_3__leaf_CLK ins_000_ DOUT_DAT VDD VSS
+ sg13g2_DFCNQD1
Xins_530_ RST clknet_3_4__leaf_CLK ins_083_ R[32] VDD VSS
+ sg13g2_DFCNQD1
Xins_531_ RST clknet_3_5__leaf_CLK ins_084_ R[33] VDD VSS
+ sg13g2_DFCNQD1
Xins_532_ RST clknet_3_1__leaf_CLK ins_085_ R[34] VDD VSS
+ sg13g2_DFCNQD1
Xins_533_ RST clknet_3_0__leaf_CLK ins_086_ R[35] VDD VSS
+ sg13g2_DFCNQD1
Xins_534_ RST clknet_3_4__leaf_CLK ins_087_ R[36] VDD VSS
+ sg13g2_DFCNQD1
Xins_535_ RST clknet_3_0__leaf_CLK ins_088_ R[37] VDD VSS
+ sg13g2_DFCNQD1
Xins_536_ RST clknet_3_0__leaf_CLK ins_089_ R[38] VDD VSS
+ sg13g2_DFCNQD1
Xins_537_ RST clknet_3_4__leaf_CLK ins_090_ R[39] VDD VSS
+ sg13g2_DFCNQD1
Xins_538_ RST clknet_3_4__leaf_CLK ins_091_ R[24] VDD VSS
+ sg13g2_DFCNQD1
Xins_539_ RST clknet_3_4__leaf_CLK ins_092_ R[25] VDD VSS
+ sg13g2_DFCNQD1
Xins_540_ RST clknet_3_1__leaf_CLK ins_093_ R[26] VDD VSS
+ sg13g2_DFCNQD1
Xins_541_ RST clknet_3_1__leaf_CLK ins_094_ R[27] VDD VSS
+ sg13g2_DFCNQD1
Xins_542_ RST clknet_3_1__leaf_CLK ins_095_ R[28] VDD VSS
+ sg13g2_DFCNQD1
Xins_543_ RST clknet_3_4__leaf_CLK ins_096_ R[29] VDD VSS
+ sg13g2_DFCNQD1
Xins_544_ RST clknet_3_1__leaf_CLK ins_097_ R[30] VDD VSS
+ sg13g2_DFCNQD1
Xins_545_ RST clknet_3_1__leaf_CLK ins_098_ R[31] VDD VSS
+ sg13g2_DFCNQD1
Xins_546_ RST clknet_3_1__leaf_CLK ins_099_ R[8] VDD VSS sg13g2_DFCNQD1
Xins_547_ RST clknet_3_5__leaf_CLK ins_100_ R[9] VDD VSS sg13g2_DFCNQD1
Xins_548_ RST clknet_3_5__leaf_CLK ins_101_ R[10] VDD VSS
+ sg13g2_DFCNQD1
Xins_549_ RST clknet_3_1__leaf_CLK ins_102_ R[11] VDD VSS
+ sg13g2_DFCNQD1
Xins_550_ RST clknet_3_0__leaf_CLK ins_103_ R[12] VDD VSS
+ sg13g2_DFCNQD1
Xins_551_ RST clknet_3_0__leaf_CLK ins_104_ R[13] VDD VSS
+ sg13g2_DFCNQD1
Xins_552_ RST clknet_3_4__leaf_CLK ins_105_ R[14] VDD VSS
+ sg13g2_DFCNQD1
Xins_553_ RST clknet_3_0__leaf_CLK ins_106_ R[15] VDD VSS
+ sg13g2_DFCNQD1
Xins_554_ RST clknet_3_6__leaf_CLK ins_107_ re VDD VSS sg13g2_DFCNQD1
Xclkbuf_0_CLK CLK VDD VSS clknet_0_CLK sg13g2_BUFFD1
Xclkbuf_3_0__f_CLK clknet_0_CLK VDD VSS clknet_3_0__leaf_CLK
+ sg13g2_BUFFD1
Xclkbuf_3_1__f_CLK clknet_0_CLK VDD VSS clknet_3_1__leaf_CLK
+ sg13g2_BUFFD1
Xclkbuf_3_2__f_CLK clknet_0_CLK VDD VSS clknet_3_2__leaf_CLK
+ sg13g2_BUFFD1
Xclkbuf_3_3__f_CLK clknet_0_CLK VDD VSS clknet_3_3__leaf_CLK
+ sg13g2_BUFFD1
Xclkbuf_3_4__f_CLK clknet_0_CLK VDD VSS clknet_3_4__leaf_CLK
+ sg13g2_BUFFD1
Xclkbuf_3_5__f_CLK clknet_0_CLK VDD VSS clknet_3_5__leaf_CLK
+ sg13g2_BUFFD1
Xclkbuf_3_6__f_CLK clknet_0_CLK VDD VSS clknet_3_6__leaf_CLK
+ sg13g2_BUFFD1
Xclkbuf_3_7__f_CLK clknet_0_CLK VDD VSS clknet_3_7__leaf_CLK
+ sg13g2_BUFFD1
Xclkload0 clknet_3_1__leaf_CLK _unconnected_0 VSS VDD sg13g2_INVD1
Xclkload1 clknet_3_2__leaf_CLK _unconnected_1 VSS VDD sg13g2_INVD1
Xclkload2 clknet_3_3__leaf_CLK _unconnected_2 VSS VDD sg13g2_INVD1
Xclkload3 clknet_3_4__leaf_CLK _unconnected_3 VSS VDD sg13g2_INVD1
Xclkload4 clknet_3_5__leaf_CLK _unconnected_4 VSS VDD sg13g2_INVD1
Xclkload5 clknet_3_6__leaf_CLK _unconnected_5 VSS VDD sg13g2_INVD1
Xclkload6 clknet_3_7__leaf_CLK _unconnected_6 VSS VDD sg13g2_INVD1
XFILLER_0_50 VDD VSS sg13g2_FILL8
XFILLER_0_58 VDD VSS sg13g2_FILL4
XFILLER_0_128 VDD VSS sg13g2_FILL8
XFILLER_0_136 VDD VSS sg13g2_FILL1
XFILLER_0_153 VDD VSS sg13g2_FILL8
XFILLER_0_161 VDD VSS sg13g2_FILL2
XFILLER_0_176 VDD VSS sg13g2_FILL1
XFILLER_0_206 VDD VSS sg13g2_FILL2
XFILLER_0_229 VDD VSS sg13g2_FILL4
XFILLER_0_275 VDD VSS sg13g2_FILL1
XFILLER_0_297 VDD VSS sg13g2_FILL4
XFILLER_0_301 VDD VSS sg13g2_FILL1
XFILLER_0_344 VDD VSS sg13g2_FILL4
XFILLER_0_348 VDD VSS sg13g2_FILL1
XFILLER_0_381 VDD VSS sg13g2_FILL4
XFILLER_0_457 VDD VSS sg13g2_FILL8
XFILLER_0_465 VDD VSS sg13g2_FILL1
XFILLER_1_0 VDD VSS sg13g2_FILL2
XFILLER_1_284 VDD VSS sg13g2_FILL4
XFILLER_1_288 VDD VSS sg13g2_FILL1
XFILLER_1_305 VDD VSS sg13g2_FILL1
XFILLER_1_335 VDD VSS sg13g2_FILL4
XFILLER_1_339 VDD VSS sg13g2_FILL2
XFILLER_1_386 VDD VSS sg13g2_FILL2
XFILLER_1_460 VDD VSS sg13g2_FILL4
XFILLER_1_464 VDD VSS sg13g2_FILL2
XFILLER_2_94 VDD VSS sg13g2_FILL4
XFILLER_2_158 VDD VSS sg13g2_FILL8
XFILLER_2_232 VDD VSS sg13g2_FILL4
XFILLER_2_236 VDD VSS sg13g2_FILL2
XFILLER_2_238 VDD VSS sg13g2_FILL1
XFILLER_2_252 VDD VSS sg13g2_FILL4
XFILLER_2_256 VDD VSS sg13g2_FILL2
XFILLER_2_364 VDD VSS sg13g2_FILL2
XFILLER_2_460 VDD VSS sg13g2_FILL4
XFILLER_2_464 VDD VSS sg13g2_FILL2
XFILLER_3_0 VDD VSS sg13g2_FILL2
XFILLER_3_162 VDD VSS sg13g2_FILL4
XFILLER_3_166 VDD VSS sg13g2_FILL2
XFILLER_3_168 VDD VSS sg13g2_FILL1
XFILLER_3_277 VDD VSS sg13g2_FILL1
XFILLER_3_305 VDD VSS sg13g2_FILL1
XFILLER_3_322 VDD VSS sg13g2_FILL4
XFILLER_3_326 VDD VSS sg13g2_FILL2
XFILLER_3_328 VDD VSS sg13g2_FILL1
XFILLER_3_355 VDD VSS sg13g2_FILL4
XFILLER_3_359 VDD VSS sg13g2_FILL2
XFILLER_3_361 VDD VSS sg13g2_FILL1
XFILLER_3_408 VDD VSS sg13g2_FILL2
XFILLER_3_410 VDD VSS sg13g2_FILL1
XFILLER_3_461 VDD VSS sg13g2_FILL4
XFILLER_3_465 VDD VSS sg13g2_FILL1
XFILLER_4_0 VDD VSS sg13g2_FILL4
XFILLER_4_4 VDD VSS sg13g2_FILL2
XFILLER_4_78 VDD VSS sg13g2_FILL4
XFILLER_4_82 VDD VSS sg13g2_FILL1
XFILLER_4_105 VDD VSS sg13g2_FILL8
XFILLER_4_113 VDD VSS sg13g2_FILL1
XFILLER_4_164 VDD VSS sg13g2_FILL8
XFILLER_4_172 VDD VSS sg13g2_FILL4
XFILLER_4_192 VDD VSS sg13g2_FILL2
XFILLER_4_207 VDD VSS sg13g2_FILL8
XFILLER_4_331 VDD VSS sg13g2_FILL2
XFILLER_4_346 VDD VSS sg13g2_FILL2
XFILLER_4_348 VDD VSS sg13g2_FILL1
XFILLER_4_449 VDD VSS sg13g2_FILL8
XFILLER_4_457 VDD VSS sg13g2_FILL8
XFILLER_4_465 VDD VSS sg13g2_FILL1
XFILLER_5_0 VDD VSS sg13g2_FILL8
XFILLER_5_8 VDD VSS sg13g2_FILL8
XFILLER_5_16 VDD VSS sg13g2_FILL1
XFILLER_5_67 VDD VSS sg13g2_FILL4
XFILLER_5_71 VDD VSS sg13g2_FILL2
XFILLER_5_123 VDD VSS sg13g2_FILL4
XFILLER_5_127 VDD VSS sg13g2_FILL2
XFILLER_5_129 VDD VSS sg13g2_FILL1
XFILLER_5_241 VDD VSS sg13g2_FILL1
XFILLER_5_264 VDD VSS sg13g2_FILL8
XFILLER_5_272 VDD VSS sg13g2_FILL4
XFILLER_5_276 VDD VSS sg13g2_FILL1
XFILLER_5_385 VDD VSS sg13g2_FILL4
XFILLER_5_389 VDD VSS sg13g2_FILL2
XFILLER_5_463 VDD VSS sg13g2_FILL2
XFILLER_5_465 VDD VSS sg13g2_FILL1
XFILLER_6_264 VDD VSS sg13g2_FILL8
XFILLER_6_272 VDD VSS sg13g2_FILL8
XFILLER_6_280 VDD VSS sg13g2_FILL2
XFILLER_6_282 VDD VSS sg13g2_FILL1
XFILLER_6_321 VDD VSS sg13g2_FILL8
XFILLER_6_329 VDD VSS sg13g2_FILL2
XFILLER_6_331 VDD VSS sg13g2_FILL1
XFILLER_6_345 VDD VSS sg13g2_FILL2
XFILLER_6_347 VDD VSS sg13g2_FILL1
XFILLER_6_383 VDD VSS sg13g2_FILL8
XFILLER_6_391 VDD VSS sg13g2_FILL1
XFILLER_6_464 VDD VSS sg13g2_FILL2
XFILLER_7_0 VDD VSS sg13g2_FILL8
XFILLER_7_8 VDD VSS sg13g2_FILL2
XFILLER_7_62 VDD VSS sg13g2_FILL4
XFILLER_7_166 VDD VSS sg13g2_FILL2
XFILLER_7_168 VDD VSS sg13g2_FILL1
XFILLER_7_182 VDD VSS sg13g2_FILL2
XFILLER_7_347 VDD VSS sg13g2_FILL8
XFILLER_7_355 VDD VSS sg13g2_FILL2
XFILLER_7_462 VDD VSS sg13g2_FILL4
XFILLER_8_0 VDD VSS sg13g2_FILL8
XFILLER_8_8 VDD VSS sg13g2_FILL2
XFILLER_8_10 VDD VSS sg13g2_FILL1
XFILLER_8_83 VDD VSS sg13g2_FILL8
XFILLER_8_91 VDD VSS sg13g2_FILL2
XFILLER_8_93 VDD VSS sg13g2_FILL1
XFILLER_8_116 VDD VSS sg13g2_FILL4
XFILLER_8_120 VDD VSS sg13g2_FILL2
XFILLER_8_122 VDD VSS sg13g2_FILL1
XFILLER_8_216 VDD VSS sg13g2_FILL4
XFILLER_8_220 VDD VSS sg13g2_FILL2
XFILLER_8_222 VDD VSS sg13g2_FILL1
XFILLER_8_245 VDD VSS sg13g2_FILL2
XFILLER_8_269 VDD VSS sg13g2_FILL8
XFILLER_8_277 VDD VSS sg13g2_FILL2
XFILLER_8_318 VDD VSS sg13g2_FILL8
XFILLER_8_326 VDD VSS sg13g2_FILL4
XFILLER_8_432 VDD VSS sg13g2_FILL8
XFILLER_8_440 VDD VSS sg13g2_FILL8
XFILLER_8_448 VDD VSS sg13g2_FILL8
XFILLER_8_456 VDD VSS sg13g2_FILL8
XFILLER_8_464 VDD VSS sg13g2_FILL2
XFILLER_9_0 VDD VSS sg13g2_FILL8
XFILLER_9_8 VDD VSS sg13g2_FILL2
XFILLER_9_60 VDD VSS sg13g2_FILL8
XFILLER_9_68 VDD VSS sg13g2_FILL4
XFILLER_9_194 VDD VSS sg13g2_FILL8
XFILLER_9_202 VDD VSS sg13g2_FILL2
XFILLER_9_204 VDD VSS sg13g2_FILL1
XFILLER_9_210 VDD VSS sg13g2_FILL8
XFILLER_9_218 VDD VSS sg13g2_FILL4
XFILLER_9_222 VDD VSS sg13g2_FILL2
XFILLER_9_246 VDD VSS sg13g2_FILL8
XFILLER_9_276 VDD VSS sg13g2_FILL4
XFILLER_9_302 VDD VSS sg13g2_FILL2
XFILLER_9_330 VDD VSS sg13g2_FILL2
XFILLER_9_345 VDD VSS sg13g2_FILL4
XFILLER_9_371 VDD VSS sg13g2_FILL8
XFILLER_9_379 VDD VSS sg13g2_FILL8
XFILLER_9_387 VDD VSS sg13g2_FILL2
XFILLER_9_461 VDD VSS sg13g2_FILL4
XFILLER_9_465 VDD VSS sg13g2_FILL1
XFILLER_10_0 VDD VSS sg13g2_FILL8
XFILLER_10_8 VDD VSS sg13g2_FILL8
XFILLER_10_132 VDD VSS sg13g2_FILL2
XFILLER_10_134 VDD VSS sg13g2_FILL1
XFILLER_10_170 VDD VSS sg13g2_FILL2
XFILLER_10_172 VDD VSS sg13g2_FILL1
XFILLER_10_178 VDD VSS sg13g2_FILL4
XFILLER_10_182 VDD VSS sg13g2_FILL2
XFILLER_10_184 VDD VSS sg13g2_FILL1
XFILLER_10_262 VDD VSS sg13g2_FILL8
XFILLER_10_270 VDD VSS sg13g2_FILL4
XFILLER_10_274 VDD VSS sg13g2_FILL2
XFILLER_10_276 VDD VSS sg13g2_FILL1
XFILLER_10_377 VDD VSS sg13g2_FILL8
XFILLER_10_385 VDD VSS sg13g2_FILL4
XFILLER_10_461 VDD VSS sg13g2_FILL4
XFILLER_10_465 VDD VSS sg13g2_FILL1
XFILLER_11_0 VDD VSS sg13g2_FILL1
XFILLER_11_51 VDD VSS sg13g2_FILL8
XFILLER_11_59 VDD VSS sg13g2_FILL8
XFILLER_11_67 VDD VSS sg13g2_FILL4
XFILLER_11_121 VDD VSS sg13g2_FILL8
XFILLER_11_129 VDD VSS sg13g2_FILL8
XFILLER_11_137 VDD VSS sg13g2_FILL2
XFILLER_11_189 VDD VSS sg13g2_FILL4
XFILLER_11_293 VDD VSS sg13g2_FILL4
XFILLER_11_297 VDD VSS sg13g2_FILL2
XFILLER_11_299 VDD VSS sg13g2_FILL1
XFILLER_11_375 VDD VSS sg13g2_FILL2
XFILLER_11_437 VDD VSS sg13g2_FILL8
XFILLER_11_445 VDD VSS sg13g2_FILL8
XFILLER_11_453 VDD VSS sg13g2_FILL8
XFILLER_11_461 VDD VSS sg13g2_FILL4
XFILLER_11_465 VDD VSS sg13g2_FILL1
XFILLER_12_0 VDD VSS sg13g2_FILL8
XFILLER_12_8 VDD VSS sg13g2_FILL8
XFILLER_12_16 VDD VSS sg13g2_FILL2
XFILLER_12_118 VDD VSS sg13g2_FILL8
XFILLER_12_198 VDD VSS sg13g2_FILL8
XFILLER_12_206 VDD VSS sg13g2_FILL8
XFILLER_12_214 VDD VSS sg13g2_FILL8
XFILLER_12_222 VDD VSS sg13g2_FILL8
XFILLER_12_230 VDD VSS sg13g2_FILL2
XFILLER_12_232 VDD VSS sg13g2_FILL1
XFILLER_12_241 VDD VSS sg13g2_FILL2
XFILLER_12_243 VDD VSS sg13g2_FILL1
XFILLER_12_266 VDD VSS sg13g2_FILL8
XFILLER_12_274 VDD VSS sg13g2_FILL8
XFILLER_12_282 VDD VSS sg13g2_FILL4
XFILLER_12_308 VDD VSS sg13g2_FILL2
XFILLER_12_310 VDD VSS sg13g2_FILL1
XFILLER_12_341 VDD VSS sg13g2_FILL1
XFILLER_12_405 VDD VSS sg13g2_FILL8
XFILLER_12_413 VDD VSS sg13g2_FILL2
XFILLER_12_415 VDD VSS sg13g2_FILL1
XFILLER_13_0 VDD VSS sg13g2_FILL8
XFILLER_13_8 VDD VSS sg13g2_FILL4
XFILLER_13_62 VDD VSS sg13g2_FILL8
XFILLER_13_70 VDD VSS sg13g2_FILL4
XFILLER_13_74 VDD VSS sg13g2_FILL1
XFILLER_13_147 VDD VSS sg13g2_FILL8
XFILLER_13_155 VDD VSS sg13g2_FILL4
XFILLER_13_159 VDD VSS sg13g2_FILL2
XFILLER_13_383 VDD VSS sg13g2_FILL8
XFILLER_13_391 VDD VSS sg13g2_FILL4
XFILLER_13_439 VDD VSS sg13g2_FILL8
XFILLER_13_447 VDD VSS sg13g2_FILL8
XFILLER_13_455 VDD VSS sg13g2_FILL8
XFILLER_13_463 VDD VSS sg13g2_FILL2
XFILLER_13_465 VDD VSS sg13g2_FILL1
XFILLER_14_0 VDD VSS sg13g2_FILL8
XFILLER_14_8 VDD VSS sg13g2_FILL4
XFILLER_14_12 VDD VSS sg13g2_FILL2
XFILLER_14_86 VDD VSS sg13g2_FILL4
XFILLER_14_184 VDD VSS sg13g2_FILL8
XFILLER_14_242 VDD VSS sg13g2_FILL8
XFILLER_14_250 VDD VSS sg13g2_FILL2
XFILLER_14_302 VDD VSS sg13g2_FILL4
XFILLER_14_314 VDD VSS sg13g2_FILL2
XFILLER_14_316 VDD VSS sg13g2_FILL1
XFILLER_14_367 VDD VSS sg13g2_FILL8
XFILLER_14_375 VDD VSS sg13g2_FILL4
XFILLER_14_379 VDD VSS sg13g2_FILL2
XFILLER_14_403 VDD VSS sg13g2_FILL8
XFILLER_14_411 VDD VSS sg13g2_FILL4
XFILLER_14_415 VDD VSS sg13g2_FILL1
XFILLER_15_0 VDD VSS sg13g2_FILL8
XFILLER_15_8 VDD VSS sg13g2_FILL4
XFILLER_15_12 VDD VSS sg13g2_FILL2
XFILLER_15_14 VDD VSS sg13g2_FILL1
XFILLER_15_37 VDD VSS sg13g2_FILL8
XFILLER_15_45 VDD VSS sg13g2_FILL8
XFILLER_15_125 VDD VSS sg13g2_FILL8
XFILLER_15_133 VDD VSS sg13g2_FILL8
XFILLER_15_141 VDD VSS sg13g2_FILL2
XFILLER_15_215 VDD VSS sg13g2_FILL8
XFILLER_15_223 VDD VSS sg13g2_FILL8
XFILLER_15_231 VDD VSS sg13g2_FILL8
XFILLER_15_239 VDD VSS sg13g2_FILL8
XFILLER_15_291 VDD VSS sg13g2_FILL4
XFILLER_15_295 VDD VSS sg13g2_FILL1
XFILLER_15_362 VDD VSS sg13g2_FILL8
XFILLER_15_370 VDD VSS sg13g2_FILL8
XFILLER_15_378 VDD VSS sg13g2_FILL2
XFILLER_15_380 VDD VSS sg13g2_FILL1
XFILLER_15_431 VDD VSS sg13g2_FILL8
XFILLER_15_439 VDD VSS sg13g2_FILL8
XFILLER_15_447 VDD VSS sg13g2_FILL8
XFILLER_15_455 VDD VSS sg13g2_FILL8
XFILLER_15_463 VDD VSS sg13g2_FILL2
XFILLER_15_465 VDD VSS sg13g2_FILL1
XFILLER_16_0 VDD VSS sg13g2_FILL8
XFILLER_16_8 VDD VSS sg13g2_FILL2
XFILLER_16_10 VDD VSS sg13g2_FILL1
XFILLER_16_61 VDD VSS sg13g2_FILL4
XFILLER_16_65 VDD VSS sg13g2_FILL2
XFILLER_16_67 VDD VSS sg13g2_FILL1
XFILLER_16_118 VDD VSS sg13g2_FILL8
XFILLER_16_126 VDD VSS sg13g2_FILL8
XFILLER_16_134 VDD VSS sg13g2_FILL4
XFILLER_16_160 VDD VSS sg13g2_FILL8
XFILLER_16_168 VDD VSS sg13g2_FILL8
XFILLER_16_176 VDD VSS sg13g2_FILL4
XFILLER_16_180 VDD VSS sg13g2_FILL1
XFILLER_16_203 VDD VSS sg13g2_FILL1
XFILLER_16_420 VDD VSS sg13g2_FILL8
XFILLER_16_428 VDD VSS sg13g2_FILL8
XFILLER_16_436 VDD VSS sg13g2_FILL8
XFILLER_16_444 VDD VSS sg13g2_FILL8
XFILLER_16_452 VDD VSS sg13g2_FILL8
XFILLER_16_460 VDD VSS sg13g2_FILL4
XFILLER_16_464 VDD VSS sg13g2_FILL2
XFILLER_17_0 VDD VSS sg13g2_FILL8
XFILLER_17_8 VDD VSS sg13g2_FILL4
XFILLER_17_62 VDD VSS sg13g2_FILL1
XFILLER_17_113 VDD VSS sg13g2_FILL2
XFILLER_17_115 VDD VSS sg13g2_FILL1
XFILLER_17_266 VDD VSS sg13g2_FILL8
XFILLER_17_274 VDD VSS sg13g2_FILL8
XFILLER_17_282 VDD VSS sg13g2_FILL8
XFILLER_17_290 VDD VSS sg13g2_FILL8
XFILLER_17_298 VDD VSS sg13g2_FILL8
XFILLER_17_306 VDD VSS sg13g2_FILL8
XFILLER_17_314 VDD VSS sg13g2_FILL8
XFILLER_17_322 VDD VSS sg13g2_FILL8
XFILLER_17_330 VDD VSS sg13g2_FILL8
XFILLER_17_338 VDD VSS sg13g2_FILL8
XFILLER_17_346 VDD VSS sg13g2_FILL8
XFILLER_17_354 VDD VSS sg13g2_FILL8
XFILLER_17_362 VDD VSS sg13g2_FILL8
XFILLER_17_370 VDD VSS sg13g2_FILL1
XFILLER_17_393 VDD VSS sg13g2_FILL2
XFILLER_17_413 VDD VSS sg13g2_FILL8
XFILLER_17_421 VDD VSS sg13g2_FILL8
XFILLER_17_429 VDD VSS sg13g2_FILL8
XFILLER_17_437 VDD VSS sg13g2_FILL8
XFILLER_17_445 VDD VSS sg13g2_FILL8
XFILLER_17_453 VDD VSS sg13g2_FILL8
XFILLER_17_461 VDD VSS sg13g2_FILL4
XFILLER_17_465 VDD VSS sg13g2_FILL1
XFILLER_18_0 VDD VSS sg13g2_FILL8
XFILLER_18_8 VDD VSS sg13g2_FILL8
XFILLER_18_16 VDD VSS sg13g2_FILL2
XFILLER_18_18 VDD VSS sg13g2_FILL1
XFILLER_18_41 VDD VSS sg13g2_FILL8
XFILLER_18_49 VDD VSS sg13g2_FILL2
XFILLER_18_51 VDD VSS sg13g2_FILL1
XFILLER_18_124 VDD VSS sg13g2_FILL8
XFILLER_18_132 VDD VSS sg13g2_FILL2
XFILLER_18_200 VDD VSS sg13g2_FILL2
XFILLER_18_267 VDD VSS sg13g2_FILL8
XFILLER_18_275 VDD VSS sg13g2_FILL8
XFILLER_18_283 VDD VSS sg13g2_FILL2
XFILLER_18_328 VDD VSS sg13g2_FILL8
XFILLER_18_386 VDD VSS sg13g2_FILL2
XFILLER_18_443 VDD VSS sg13g2_FILL8
XFILLER_18_451 VDD VSS sg13g2_FILL8
XFILLER_18_459 VDD VSS sg13g2_FILL4
XFILLER_18_463 VDD VSS sg13g2_FILL2
XFILLER_18_465 VDD VSS sg13g2_FILL1
XFILLER_19_0 VDD VSS sg13g2_FILL8
XFILLER_19_8 VDD VSS sg13g2_FILL4
XFILLER_19_12 VDD VSS sg13g2_FILL2
XFILLER_19_14 VDD VSS sg13g2_FILL1
XFILLER_19_37 VDD VSS sg13g2_FILL8
XFILLER_19_45 VDD VSS sg13g2_FILL8
XFILLER_19_53 VDD VSS sg13g2_FILL4
XFILLER_19_57 VDD VSS sg13g2_FILL1
XFILLER_19_93 VDD VSS sg13g2_FILL8
XFILLER_19_101 VDD VSS sg13g2_FILL2
XFILLER_19_103 VDD VSS sg13g2_FILL1
XFILLER_19_148 VDD VSS sg13g2_FILL4
XFILLER_19_152 VDD VSS sg13g2_FILL2
XFILLER_19_388 VDD VSS sg13g2_FILL4
XFILLER_19_450 VDD VSS sg13g2_FILL8
XFILLER_19_458 VDD VSS sg13g2_FILL8
XFILLER_20_0 VDD VSS sg13g2_FILL8
XFILLER_20_8 VDD VSS sg13g2_FILL8
XFILLER_20_16 VDD VSS sg13g2_FILL8
XFILLER_20_24 VDD VSS sg13g2_FILL8
XFILLER_20_32 VDD VSS sg13g2_FILL8
XFILLER_20_40 VDD VSS sg13g2_FILL8
XFILLER_20_48 VDD VSS sg13g2_FILL8
XFILLER_20_56 VDD VSS sg13g2_FILL8
XFILLER_20_64 VDD VSS sg13g2_FILL8
XFILLER_20_72 VDD VSS sg13g2_FILL8
XFILLER_20_80 VDD VSS sg13g2_FILL8
XFILLER_20_88 VDD VSS sg13g2_FILL8
XFILLER_20_96 VDD VSS sg13g2_FILL8
XFILLER_20_104 VDD VSS sg13g2_FILL4
XFILLER_20_108 VDD VSS sg13g2_FILL1
XFILLER_20_167 VDD VSS sg13g2_FILL2
XFILLER_20_191 VDD VSS sg13g2_FILL8
XFILLER_20_199 VDD VSS sg13g2_FILL2
XFILLER_20_251 VDD VSS sg13g2_FILL8
XFILLER_20_259 VDD VSS sg13g2_FILL8
XFILLER_20_438 VDD VSS sg13g2_FILL8
XFILLER_20_446 VDD VSS sg13g2_FILL8
XFILLER_20_454 VDD VSS sg13g2_FILL8
XFILLER_20_462 VDD VSS sg13g2_FILL4
XFILLER_21_0 VDD VSS sg13g2_FILL8
XFILLER_21_8 VDD VSS sg13g2_FILL8
XFILLER_21_16 VDD VSS sg13g2_FILL8
XFILLER_21_24 VDD VSS sg13g2_FILL8
XFILLER_21_32 VDD VSS sg13g2_FILL8
XFILLER_21_40 VDD VSS sg13g2_FILL8
XFILLER_21_48 VDD VSS sg13g2_FILL8
XFILLER_21_56 VDD VSS sg13g2_FILL8
XFILLER_21_64 VDD VSS sg13g2_FILL8
XFILLER_21_72 VDD VSS sg13g2_FILL8
XFILLER_21_80 VDD VSS sg13g2_FILL8
XFILLER_21_88 VDD VSS sg13g2_FILL8
XFILLER_21_96 VDD VSS sg13g2_FILL8
XFILLER_21_180 VDD VSS sg13g2_FILL8
XFILLER_21_188 VDD VSS sg13g2_FILL4
XFILLER_21_205 VDD VSS sg13g2_FILL2
XFILLER_21_207 VDD VSS sg13g2_FILL1
XFILLER_21_244 VDD VSS sg13g2_FILL8
XFILLER_21_252 VDD VSS sg13g2_FILL8
XFILLER_21_260 VDD VSS sg13g2_FILL2
XFILLER_21_262 VDD VSS sg13g2_FILL1
XFILLER_21_276 VDD VSS sg13g2_FILL4
XFILLER_21_280 VDD VSS sg13g2_FILL2
XFILLER_21_282 VDD VSS sg13g2_FILL1
XFILLER_21_291 VDD VSS sg13g2_FILL8
XFILLER_21_299 VDD VSS sg13g2_FILL8
XFILLER_21_307 VDD VSS sg13g2_FILL1
XFILLER_21_359 VDD VSS sg13g2_FILL1
XFILLER_21_389 VDD VSS sg13g2_FILL2
XFILLER_21_441 VDD VSS sg13g2_FILL8
XFILLER_21_449 VDD VSS sg13g2_FILL8
XFILLER_21_457 VDD VSS sg13g2_FILL8
XFILLER_21_465 VDD VSS sg13g2_FILL1
XFILLER_22_0 VDD VSS sg13g2_FILL8
XFILLER_22_8 VDD VSS sg13g2_FILL8
XFILLER_22_16 VDD VSS sg13g2_FILL8
XFILLER_22_24 VDD VSS sg13g2_FILL8
XFILLER_22_32 VDD VSS sg13g2_FILL8
XFILLER_22_40 VDD VSS sg13g2_FILL8
XFILLER_22_48 VDD VSS sg13g2_FILL8
XFILLER_22_56 VDD VSS sg13g2_FILL8
XFILLER_22_64 VDD VSS sg13g2_FILL8
XFILLER_22_72 VDD VSS sg13g2_FILL8
XFILLER_22_80 VDD VSS sg13g2_FILL8
XFILLER_22_88 VDD VSS sg13g2_FILL8
XFILLER_22_96 VDD VSS sg13g2_FILL8
XFILLER_22_104 VDD VSS sg13g2_FILL4
XFILLER_22_108 VDD VSS sg13g2_FILL2
XFILLER_22_110 VDD VSS sg13g2_FILL1
XFILLER_22_182 VDD VSS sg13g2_FILL2
XFILLER_22_208 VDD VSS sg13g2_FILL2
XFILLER_22_210 VDD VSS sg13g2_FILL1
XFILLER_22_311 VDD VSS sg13g2_FILL4
XFILLER_22_315 VDD VSS sg13g2_FILL2
XFILLER_22_367 VDD VSS sg13g2_FILL1
XFILLER_22_418 VDD VSS sg13g2_FILL8
XFILLER_22_426 VDD VSS sg13g2_FILL8
XFILLER_22_434 VDD VSS sg13g2_FILL8
XFILLER_22_442 VDD VSS sg13g2_FILL8
XFILLER_22_450 VDD VSS sg13g2_FILL8
XFILLER_22_458 VDD VSS sg13g2_FILL8
XFILLER_23_0 VDD VSS sg13g2_FILL8
XFILLER_23_8 VDD VSS sg13g2_FILL8
XFILLER_23_16 VDD VSS sg13g2_FILL8
XFILLER_23_24 VDD VSS sg13g2_FILL8
XFILLER_23_32 VDD VSS sg13g2_FILL8
XFILLER_23_40 VDD VSS sg13g2_FILL8
XFILLER_23_48 VDD VSS sg13g2_FILL8
XFILLER_23_56 VDD VSS sg13g2_FILL8
XFILLER_23_64 VDD VSS sg13g2_FILL8
XFILLER_23_72 VDD VSS sg13g2_FILL8
XFILLER_23_80 VDD VSS sg13g2_FILL8
XFILLER_23_88 VDD VSS sg13g2_FILL8
XFILLER_23_96 VDD VSS sg13g2_FILL8
XFILLER_23_104 VDD VSS sg13g2_FILL8
XFILLER_23_112 VDD VSS sg13g2_FILL1
XFILLER_23_423 VDD VSS sg13g2_FILL8
XFILLER_23_431 VDD VSS sg13g2_FILL8
XFILLER_23_439 VDD VSS sg13g2_FILL8
XFILLER_23_447 VDD VSS sg13g2_FILL8
XFILLER_23_455 VDD VSS sg13g2_FILL8
XFILLER_23_463 VDD VSS sg13g2_FILL2
XFILLER_23_465 VDD VSS sg13g2_FILL1
XFILLER_24_0 VDD VSS sg13g2_FILL8
XFILLER_24_8 VDD VSS sg13g2_FILL8
XFILLER_24_16 VDD VSS sg13g2_FILL8
XFILLER_24_24 VDD VSS sg13g2_FILL8
XFILLER_24_32 VDD VSS sg13g2_FILL8
XFILLER_24_40 VDD VSS sg13g2_FILL8
XFILLER_24_48 VDD VSS sg13g2_FILL8
XFILLER_24_56 VDD VSS sg13g2_FILL8
XFILLER_24_64 VDD VSS sg13g2_FILL8
XFILLER_24_72 VDD VSS sg13g2_FILL8
XFILLER_24_80 VDD VSS sg13g2_FILL8
XFILLER_24_88 VDD VSS sg13g2_FILL8
XFILLER_24_96 VDD VSS sg13g2_FILL8
XFILLER_24_104 VDD VSS sg13g2_FILL8
XFILLER_24_112 VDD VSS sg13g2_FILL8
XFILLER_24_120 VDD VSS sg13g2_FILL1
XFILLER_24_171 VDD VSS sg13g2_FILL8
XFILLER_24_179 VDD VSS sg13g2_FILL2
XFILLER_24_244 VDD VSS sg13g2_FILL8
XFILLER_24_252 VDD VSS sg13g2_FILL8
XFILLER_24_260 VDD VSS sg13g2_FILL8
XFILLER_24_268 VDD VSS sg13g2_FILL8
XFILLER_24_276 VDD VSS sg13g2_FILL2
XFILLER_24_291 VDD VSS sg13g2_FILL8
XFILLER_24_320 VDD VSS sg13g2_FILL4
XFILLER_24_324 VDD VSS sg13g2_FILL1
XFILLER_24_338 VDD VSS sg13g2_FILL8
XFILLER_24_346 VDD VSS sg13g2_FILL2
XFILLER_24_369 VDD VSS sg13g2_FILL8
XFILLER_24_377 VDD VSS sg13g2_FILL8
XFILLER_24_393 VDD VSS sg13g2_FILL8
XFILLER_24_401 VDD VSS sg13g2_FILL8
XFILLER_24_409 VDD VSS sg13g2_FILL8
XFILLER_24_417 VDD VSS sg13g2_FILL8
XFILLER_24_425 VDD VSS sg13g2_FILL8
XFILLER_24_433 VDD VSS sg13g2_FILL8
XFILLER_24_441 VDD VSS sg13g2_FILL8
XFILLER_24_449 VDD VSS sg13g2_FILL8
XFILLER_24_457 VDD VSS sg13g2_FILL8
XFILLER_24_465 VDD VSS sg13g2_FILL1
.ENDS SPI
* CDL Netlist generated by OpenROAD

*.BUSDELIMITER [

.SUBCKT asicone_202508 AVDD VDD VDDIO VSS VSSIO pad_adc_clk_pad
+ pad_adc_go_pad pad_adc_result_0_pad pad_adc_result_1_pad pad_adc_result_2_pad
+ pad_adc_result_3_pad pad_adc_result_4_pad pad_adc_rst_pad
+ pad_adc_sample_pad pad_adc_valid_pad pad_adc_vin_pad pad_adc_vip_pad
+ pad_adc_vrefn_pad pad_adc_vrefp_pad pad_cs_pad pad_miso_pad
+ pad_mosi_pad pad_sclk_pad
XCORNER_1 VDDIO VSSIO VDD VSS VSS sg13g2_Corner
XCORNER_2 VDDIO VSSIO VDD VSS VSS sg13g2_Corner
XCORNER_3 VDDIO VSSIO VDD VSS VSS sg13g2_Corner
XCORNER_4 VDDIO VSSIO VDD VSS VSS sg13g2_Corner
XFILLER_0 VDDIO VSSIO VDD VSS VSS sg13g2_Filler4000
XFILLER_1 VDDIO VSSIO VDD VSS VSS sg13g2_Filler200
XFILLER_2 VDDIO VSSIO VDD VSS VSS sg13g2_Filler4000
XFILLER_3 VDDIO VSSIO VDD VSS VSS sg13g2_Filler200
XFILLER_4 VDDIO VSSIO VDD VSS VSS sg13g2_Filler4000
XFILLER_5 VDDIO VSSIO VDD VSS VSS sg13g2_Filler200
XFILLER_6 VDDIO VSSIO VDD VSS VSS sg13g2_Filler4000
XFILLER_7 VDDIO VSSIO VDD VSS VSS sg13g2_Filler200
Xadc AVDD pad_adc_clk_p2c pad_adc_go_p2c pad_adc_result_0_c2p
+ pad_adc_result_1_c2p pad_adc_result_2_c2p pad_adc_result_3_c2p
+ pad_adc_result_4_c2p pad_adc_rst_p2c pad_adc_sample_c2p pad_adc_valid_c2p
+ VDD pad_adc_vin_padres pad_adc_vip_padres pad_adc_vrefp_padres
+ pad_adc_vrefn_padres VSS SARADC
Xbd_pad_adc_avdd sg13g2_bpd70
Xbd_pad_adc_clk sg13g2_bpd70
Xbd_pad_adc_go sg13g2_bpd70
Xbd_pad_adc_result_0 sg13g2_bpd70
Xbd_pad_adc_result_1 sg13g2_bpd70
Xbd_pad_adc_result_2 sg13g2_bpd70
Xbd_pad_adc_result_3 sg13g2_bpd70
Xbd_pad_adc_result_4 sg13g2_bpd70
Xbd_pad_adc_rst sg13g2_bpd70
Xbd_pad_adc_sample sg13g2_bpd70
Xbd_pad_adc_valid sg13g2_bpd70
Xbd_pad_adc_vin sg13g2_bpd70
Xbd_pad_adc_vip sg13g2_bpd70
Xbd_pad_adc_vrefn sg13g2_bpd70
Xbd_pad_adc_vrefp sg13g2_bpd70
Xbd_pad_adc_vss sg13g2_bpd70
Xbd_pad_cs sg13g2_bpd70
Xbd_pad_dum_1 sg13g2_bpd70
Xbd_pad_dum_10 sg13g2_bpd70
Xbd_pad_dum_11 sg13g2_bpd70
Xbd_pad_dum_12 sg13g2_bpd70
Xbd_pad_dum_13 sg13g2_bpd70
Xbd_pad_dum_14 sg13g2_bpd70
Xbd_pad_dum_2 sg13g2_bpd70
Xbd_pad_dum_3 sg13g2_bpd70
Xbd_pad_dum_4 sg13g2_bpd70
Xbd_pad_dum_5 sg13g2_bpd70
Xbd_pad_dum_6 sg13g2_bpd70
Xbd_pad_dum_7 sg13g2_bpd70
Xbd_pad_dum_8 sg13g2_bpd70
Xbd_pad_dum_9 sg13g2_bpd70
Xbd_pad_miso sg13g2_bpd70
Xbd_pad_mosi sg13g2_bpd70
Xbd_pad_sclk sg13g2_bpd70
Xbd_vdd_north_0 sg13g2_bpd70
Xbd_vddpst_north_0 sg13g2_bpd70
Xbd_vss_north_0 sg13g2_bpd70
Xbd_vsspst_north_0 sg13g2_bpd70
Xbuf_spi_32 R[0] VDD VSS RD[32] sg13g2_BUFFD1
Xbuf_spi_33 R[1] VDD VSS RD[33] sg13g2_BUFFD1
Xbuf_spi_34 R[2] VDD VSS RD[34] sg13g2_BUFFD1
Xbuf_spi_35 R[3] VDD VSS RD[35] sg13g2_BUFFD1
Xbuf_spi_36 R[4] VDD VSS RD[36] sg13g2_BUFFD1
Xbuf_spi_37 R[5] VDD VSS RD[37] sg13g2_BUFFD1
Xbuf_spi_38 R[6] VDD VSS RD[38] sg13g2_BUFFD1
Xbuf_spi_39 R[7] VDD VSS RD[39] sg13g2_BUFFD1
Xbuf_spi_40 R[8] VDD VSS RD[40] sg13g2_BUFFD1
Xbuf_spi_41 R[9] VDD VSS RD[41] sg13g2_BUFFD1
Xbuf_spi_42 R[10] VDD VSS RD[42] sg13g2_BUFFD1
Xbuf_spi_43 R[11] VDD VSS RD[43] sg13g2_BUFFD1
Xbuf_spi_44 R[12] VDD VSS RD[44] sg13g2_BUFFD1
Xbuf_spi_45 R[13] VDD VSS RD[45] sg13g2_BUFFD1
Xbuf_spi_46 R[14] VDD VSS RD[46] sg13g2_BUFFD1
Xbuf_spi_47 R[15] VDD VSS RD[47] sg13g2_BUFFD1
Xpad_adc_avdd VDDIO VSSIO AVDD pad_adc_avdd_padres VDD VSS
+ VSS sg13g2_IOPadAnalog
Xpad_adc_clk VDDIO VSSIO pad_adc_clk_p2c pad_adc_clk_pad VDD
+ VSS VSS sg13g2_IOPadIn
Xpad_adc_go VDDIO VSSIO pad_adc_go_p2c pad_adc_go_pad VDD
+ VSS VSS sg13g2_IOPadIn
Xpad_adc_result_0 pad_adc_result_0_c2p VDDIO VSSIO pad_adc_result_0_pad
+ VDD VSS VSS sg13g2_IOPadOut16mA
Xpad_adc_result_1 pad_adc_result_1_c2p VDDIO VSSIO pad_adc_result_1_pad
+ VDD VSS VSS sg13g2_IOPadOut16mA
Xpad_adc_result_2 pad_adc_result_2_c2p VDDIO VSSIO pad_adc_result_2_pad
+ VDD VSS VSS sg13g2_IOPadOut16mA
Xpad_adc_result_3 pad_adc_result_3_c2p VDDIO VSSIO pad_adc_result_3_pad
+ VDD VSS VSS sg13g2_IOPadOut16mA
Xpad_adc_result_4 pad_adc_result_4_c2p VDDIO VSSIO pad_adc_result_4_pad
+ VDD VSS VSS sg13g2_IOPadOut16mA
Xpad_adc_rst VDDIO VSSIO pad_adc_rst_p2c pad_adc_rst_pad VDD
+ VSS VSS sg13g2_IOPadIn
Xpad_adc_sample pad_adc_sample_c2p VDDIO VSSIO pad_adc_sample_pad
+ VDD VSS VSS sg13g2_IOPadOut16mA
Xpad_adc_valid pad_adc_valid_c2p VDDIO VSSIO pad_adc_valid_pad
+ VDD VSS VSS sg13g2_IOPadOut16mA
Xpad_adc_vin VDDIO VSSIO pad_adc_vin_pad pad_adc_vin_padres
+ VDD VSS VSS sg13g2_IOPadAnalog
Xpad_adc_vip VDDIO VSSIO pad_adc_vip_pad pad_adc_vip_padres
+ VDD VSS VSS sg13g2_IOPadAnalog
Xpad_adc_vrefn VDDIO VSSIO pad_adc_vrefn_pad pad_adc_vrefn_padres
+ VDD VSS VSS sg13g2_IOPadAnalog
Xpad_adc_vrefp VDDIO VSSIO pad_adc_vrefp_pad pad_adc_vrefp_padres
+ VDD VSS VSS sg13g2_IOPadAnalog
Xpad_adc_vss VDDIO VSSIO VDD VSS VSS sg13g2_IOPadVssExt
Xpad_cs VDDIO VSSIO pad_cs_p2c pad_cs_pad VDD VSS VSS sg13g2_IOPadIn
Xpad_dum_1 VDDIO VSSIO _unconnected_0 _unconnected_1 VDD VSS
+ VSS sg13g2_IOPadAnalog
Xpad_dum_10 VDDIO VSSIO _unconnected_2 _unconnected_3 VDD
+ VSS VSS sg13g2_IOPadAnalog
Xpad_dum_11 VDDIO VSSIO _unconnected_4 _unconnected_5 VDD
+ VSS VSS sg13g2_IOPadAnalog
Xpad_dum_12 VDDIO VSSIO _unconnected_6 _unconnected_7 VDD
+ VSS VSS sg13g2_IOPadAnalog
Xpad_dum_13 VDDIO VSSIO _unconnected_8 _unconnected_9 VDD
+ VSS VSS sg13g2_IOPadAnalog
Xpad_dum_14 VDDIO VSSIO _unconnected_10 _unconnected_11 VDD
+ VSS VSS sg13g2_IOPadAnalog
Xpad_dum_2 VDDIO VSSIO _unconnected_12 _unconnected_13 VDD
+ VSS VSS sg13g2_IOPadAnalog
Xpad_dum_3 VDDIO VSSIO _unconnected_14 _unconnected_15 VDD
+ VSS VSS sg13g2_IOPadAnalog
Xpad_dum_4 VDDIO VSSIO _unconnected_16 _unconnected_17 VDD
+ VSS VSS sg13g2_IOPadAnalog
Xpad_dum_5 VDDIO VSSIO _unconnected_18 _unconnected_19 VDD
+ VSS VSS sg13g2_IOPadAnalog
Xpad_dum_6 VDDIO VSSIO _unconnected_20 _unconnected_21 VDD
+ VSS VSS sg13g2_IOPadAnalog
Xpad_dum_7 VDDIO VSSIO _unconnected_22 _unconnected_23 VDD
+ VSS VSS sg13g2_IOPadAnalog
Xpad_dum_8 VDDIO VSSIO _unconnected_24 _unconnected_25 VDD
+ VSS VSS sg13g2_IOPadAnalog
Xpad_dum_9 VDDIO VSSIO _unconnected_26 _unconnected_27 VDD
+ VSS VSS sg13g2_IOPadAnalog
Xpad_miso pad_miso_c2p VDDIO VSSIO pad_miso_pad VDD VSS VSS
+ sg13g2_IOPadOut16mA
Xpad_mosi VDDIO VSSIO pad_mosi_p2c pad_mosi_pad VDD VSS VSS
+ sg13g2_IOPadIn
Xpad_sclk VDDIO VSSIO pad_sclk_p2c pad_sclk_pad VDD VSS VSS
+ sg13g2_IOPadIn
Xpad_vdd_north_0 VDDIO VSSIO VDD VSS VSS sg13g2_IOPadVddExt
Xpad_vddpst_north_0 VDDIO VSSIO VDD VSS VSS sg13g2_IOPadIOVdd
Xpad_vss_north_0 VDDIO VSSIO VDD VSS VSS sg13g2_IOPadVssExt
Xpad_vsspst_north_0 VDDIO VSSIO VDD VSS VSS sg13g2_IOPadIOVss
Xspi pad_cs_p2c pad_sclk_p2c pad_mosi_p2c pad_miso_c2p _unconnected_28
+ RD[0] RD[10] RD[11] RD[12] RD[13] RD[14] RD[15] RD[16] RD[17]
+ RD[18] RD[19] RD[1] RD[20] RD[21] RD[22] RD[23] RD[24] RD[25]
+ RD[26] RD[27] RD[28] RD[29] RD[2] RD[30] RD[31] RD[32] RD[33]
+ RD[34] RD[35] RD[36] RD[37] RD[38] RD[39] RD[3] RD[40] RD[41]
+ RD[42] RD[43] RD[44] RD[45] RD[46] RD[47] RD[4] RD[5] RD[6]
+ RD[7] RD[8] RD[9] pad_adc_rst_p2c R[0] R[10] R[11] R[12] R[13]
+ R[14] R[15] R[16] R[17] R[18] R[19] R[1] R[20] R[21] R[22]
+ R[23] R[24] R[25] R[26] R[27] R[28] R[29] R[2] R[30] R[31]
+ R[32] R[33] R[34] R[35] R[36] R[37] R[38] R[39] R[3] R[40]
+ R[41] R[42] R[43] R[44] R[45] R[46] R[47] R[48] R[49] R[4]
+ R[50] R[51] R[52] R[53] R[54] R[55] R[56] R[57] R[58] R[59]
+ R[5] R[60] R[61] R[62] R[63] R[6] R[7] R[8] R[9] VSS VDD SPI
Xspi_adc_result_0 RESULT[0] VDD VSS RD[0] sg13g2_BUFFD1
Xspi_adc_result_1 RESULT[1] VDD VSS RD[1] sg13g2_BUFFD1
Xspi_adc_result_2 RESULT[2] VDD VSS RD[2] sg13g2_BUFFD1
Xspi_adc_result_3 RESULT[3] VDD VSS RD[3] sg13g2_BUFFD1
Xspi_adc_result_4 RESULT[4] VDD VSS RD[4] sg13g2_BUFFD1
Xspi_adc_sample pad_adc_sample_c2p VDD VSS RD[9] sg13g2_BUFFD1
Xspi_adc_valid pad_adc_valid_c2p VDD VSS RD[8] sg13g2_BUFFD1
Xtie_spi_0 VDD VSS RD[5] sg13g2_TIEL
Xtie_spi_1 VDD VSS RD[6] sg13g2_TIEL
Xtie_spi_10 VDD VSS RD[10] sg13g2_TIEL
Xtie_spi_11 VDD VSS RD[11] sg13g2_TIEL
Xtie_spi_12 VDD VSS RD[12] sg13g2_TIEL
Xtie_spi_13 VDD VSS RD[13] sg13g2_TIEL
Xtie_spi_14 VDD VSS RD[14] sg13g2_TIEL
Xtie_spi_15 VDD VSS RD[15] sg13g2_TIEL
Xtie_spi_16 VDD VSS RD[16] sg13g2_TIEL
Xtie_spi_17 VDD VSS RD[17] sg13g2_TIEH
Xtie_spi_18 VDD VSS RD[18] sg13g2_TIEL
Xtie_spi_19 VDD VSS RD[19] sg13g2_TIEH
Xtie_spi_2 VDD VSS RD[7] sg13g2_TIEL
Xtie_spi_20 VDD VSS RD[20] sg13g2_TIEL
Xtie_spi_21 VDD VSS RD[21] sg13g2_TIEH
Xtie_spi_22 VDD VSS RD[22] sg13g2_TIEL
Xtie_spi_23 VDD VSS RD[23] sg13g2_TIEH
Xtie_spi_24 VDD VSS RD[24] sg13g2_TIEH
Xtie_spi_25 VDD VSS RD[25] sg13g2_TIEL
Xtie_spi_26 VDD VSS RD[26] sg13g2_TIEH
Xtie_spi_27 VDD VSS RD[27] sg13g2_TIEL
Xtie_spi_28 VDD VSS RD[28] sg13g2_TIEH
Xtie_spi_29 VDD VSS RD[29] sg13g2_TIEL
Xtie_spi_30 VDD VSS RD[30] sg13g2_TIEH
Xtie_spi_31 VDD VSS RD[31] sg13g2_TIEL
XANTENNA_1 pad_adc_sample_c2p VDD VSS sg13g2_ANTENNA
XANTENNA_2 pad_adc_sample_c2p VDD VSS sg13g2_ANTENNA
XANTENNA_3 pad_adc_valid_c2p VDD VSS sg13g2_ANTENNA
XANTENNA_4 pad_adc_valid_c2p VDD VSS sg13g2_ANTENNA
XSTDFILL0_0 VDD VSS sg13g2_FILL8
XSTDFILL0_8 VDD VSS sg13g2_FILL8
XSTDFILL0_16 VDD VSS sg13g2_FILL8
XSTDFILL0_24 VDD VSS sg13g2_FILL8
XSTDFILL0_32 VDD VSS sg13g2_FILL8
XSTDFILL0_40 VDD VSS sg13g2_FILL8
XSTDFILL0_48 VDD VSS sg13g2_FILL8
XSTDFILL0_56 VDD VSS sg13g2_FILL8
XSTDFILL0_64 VDD VSS sg13g2_FILL8
XSTDFILL0_72 VDD VSS sg13g2_FILL8
XSTDFILL0_80 VDD VSS sg13g2_FILL8
XSTDFILL0_88 VDD VSS sg13g2_FILL8
XSTDFILL0_96 VDD VSS sg13g2_FILL8
XSTDFILL0_104 VDD VSS sg13g2_FILL1
XSTDFILL0_1880 VDD VSS sg13g2_FILL8
XSTDFILL0_1888 VDD VSS sg13g2_FILL8
XSTDFILL0_1896 VDD VSS sg13g2_FILL8
XSTDFILL0_1904 VDD VSS sg13g2_FILL8
XSTDFILL0_1912 VDD VSS sg13g2_FILL8
XSTDFILL0_1920 VDD VSS sg13g2_FILL8
XSTDFILL0_1928 VDD VSS sg13g2_FILL8
XSTDFILL0_1936 VDD VSS sg13g2_FILL8
XSTDFILL0_1944 VDD VSS sg13g2_FILL8
XSTDFILL0_1952 VDD VSS sg13g2_FILL8
XSTDFILL0_1960 VDD VSS sg13g2_FILL8
XSTDFILL0_1968 VDD VSS sg13g2_FILL8
XSTDFILL0_1976 VDD VSS sg13g2_FILL8
XSTDFILL0_1984 VDD VSS sg13g2_FILL8
XSTDFILL0_1992 VDD VSS sg13g2_FILL8
XSTDFILL0_2000 VDD VSS sg13g2_FILL8
XSTDFILL0_2008 VDD VSS sg13g2_FILL8
XSTDFILL0_2016 VDD VSS sg13g2_FILL8
XSTDFILL0_2024 VDD VSS sg13g2_FILL8
XSTDFILL0_2032 VDD VSS sg13g2_FILL8
XSTDFILL0_2040 VDD VSS sg13g2_FILL8
XSTDFILL0_2048 VDD VSS sg13g2_FILL8
XSTDFILL0_2056 VDD VSS sg13g2_FILL8
XSTDFILL0_2064 VDD VSS sg13g2_FILL8
XSTDFILL0_2072 VDD VSS sg13g2_FILL8
XSTDFILL0_2080 VDD VSS sg13g2_FILL8
XSTDFILL0_2088 VDD VSS sg13g2_FILL8
XSTDFILL0_2096 VDD VSS sg13g2_FILL8
XSTDFILL0_2104 VDD VSS sg13g2_FILL8
XSTDFILL0_2112 VDD VSS sg13g2_FILL8
XSTDFILL0_2120 VDD VSS sg13g2_FILL8
XSTDFILL0_2128 VDD VSS sg13g2_FILL8
XSTDFILL0_2136 VDD VSS sg13g2_FILL8
XSTDFILL0_2144 VDD VSS sg13g2_FILL8
XSTDFILL0_2152 VDD VSS sg13g2_FILL8
XSTDFILL0_2160 VDD VSS sg13g2_FILL8
XSTDFILL0_2168 VDD VSS sg13g2_FILL4
XSTDFILL1_0 VDD VSS sg13g2_FILL8
XSTDFILL1_8 VDD VSS sg13g2_FILL8
XSTDFILL1_16 VDD VSS sg13g2_FILL8
XSTDFILL1_24 VDD VSS sg13g2_FILL8
XSTDFILL1_32 VDD VSS sg13g2_FILL8
XSTDFILL1_40 VDD VSS sg13g2_FILL8
XSTDFILL1_48 VDD VSS sg13g2_FILL8
XSTDFILL1_56 VDD VSS sg13g2_FILL8
XSTDFILL1_64 VDD VSS sg13g2_FILL8
XSTDFILL1_72 VDD VSS sg13g2_FILL8
XSTDFILL1_80 VDD VSS sg13g2_FILL8
XSTDFILL1_88 VDD VSS sg13g2_FILL8
XSTDFILL1_96 VDD VSS sg13g2_FILL8
XSTDFILL1_104 VDD VSS sg13g2_FILL1
XSTDFILL1_1880 VDD VSS sg13g2_FILL8
XSTDFILL1_1888 VDD VSS sg13g2_FILL8
XSTDFILL1_1896 VDD VSS sg13g2_FILL8
XSTDFILL1_1904 VDD VSS sg13g2_FILL8
XSTDFILL1_1912 VDD VSS sg13g2_FILL8
XSTDFILL1_1920 VDD VSS sg13g2_FILL8
XSTDFILL1_1928 VDD VSS sg13g2_FILL8
XSTDFILL1_1936 VDD VSS sg13g2_FILL8
XSTDFILL1_1944 VDD VSS sg13g2_FILL8
XSTDFILL1_1952 VDD VSS sg13g2_FILL8
XSTDFILL1_1960 VDD VSS sg13g2_FILL8
XSTDFILL1_1968 VDD VSS sg13g2_FILL8
XSTDFILL1_1976 VDD VSS sg13g2_FILL8
XSTDFILL1_1984 VDD VSS sg13g2_FILL8
XSTDFILL1_1992 VDD VSS sg13g2_FILL8
XSTDFILL1_2000 VDD VSS sg13g2_FILL8
XSTDFILL1_2008 VDD VSS sg13g2_FILL8
XSTDFILL1_2016 VDD VSS sg13g2_FILL8
XSTDFILL1_2024 VDD VSS sg13g2_FILL8
XSTDFILL1_2032 VDD VSS sg13g2_FILL8
XSTDFILL1_2040 VDD VSS sg13g2_FILL8
XSTDFILL1_2048 VDD VSS sg13g2_FILL8
XSTDFILL1_2056 VDD VSS sg13g2_FILL8
XSTDFILL1_2064 VDD VSS sg13g2_FILL8
XSTDFILL1_2072 VDD VSS sg13g2_FILL8
XSTDFILL1_2080 VDD VSS sg13g2_FILL8
XSTDFILL1_2088 VDD VSS sg13g2_FILL8
XSTDFILL1_2096 VDD VSS sg13g2_FILL8
XSTDFILL1_2104 VDD VSS sg13g2_FILL8
XSTDFILL1_2112 VDD VSS sg13g2_FILL8
XSTDFILL1_2120 VDD VSS sg13g2_FILL8
XSTDFILL1_2128 VDD VSS sg13g2_FILL8
XSTDFILL1_2136 VDD VSS sg13g2_FILL8
XSTDFILL1_2144 VDD VSS sg13g2_FILL8
XSTDFILL1_2152 VDD VSS sg13g2_FILL8
XSTDFILL1_2160 VDD VSS sg13g2_FILL8
XSTDFILL1_2168 VDD VSS sg13g2_FILL4
XSTDFILL2_0 VDD VSS sg13g2_FILL8
XSTDFILL2_8 VDD VSS sg13g2_FILL8
XSTDFILL2_16 VDD VSS sg13g2_FILL8
XSTDFILL2_24 VDD VSS sg13g2_FILL8
XSTDFILL2_32 VDD VSS sg13g2_FILL8
XSTDFILL2_40 VDD VSS sg13g2_FILL8
XSTDFILL2_48 VDD VSS sg13g2_FILL8
XSTDFILL2_56 VDD VSS sg13g2_FILL8
XSTDFILL2_64 VDD VSS sg13g2_FILL8
XSTDFILL2_72 VDD VSS sg13g2_FILL8
XSTDFILL2_80 VDD VSS sg13g2_FILL8
XSTDFILL2_88 VDD VSS sg13g2_FILL8
XSTDFILL2_96 VDD VSS sg13g2_FILL8
XSTDFILL2_104 VDD VSS sg13g2_FILL1
XSTDFILL2_1880 VDD VSS sg13g2_FILL8
XSTDFILL2_1888 VDD VSS sg13g2_FILL8
XSTDFILL2_1896 VDD VSS sg13g2_FILL8
XSTDFILL2_1904 VDD VSS sg13g2_FILL8
XSTDFILL2_1912 VDD VSS sg13g2_FILL8
XSTDFILL2_1920 VDD VSS sg13g2_FILL8
XSTDFILL2_1928 VDD VSS sg13g2_FILL8
XSTDFILL2_1936 VDD VSS sg13g2_FILL8
XSTDFILL2_1944 VDD VSS sg13g2_FILL8
XSTDFILL2_1952 VDD VSS sg13g2_FILL8
XSTDFILL2_1960 VDD VSS sg13g2_FILL8
XSTDFILL2_1968 VDD VSS sg13g2_FILL8
XSTDFILL2_1976 VDD VSS sg13g2_FILL8
XSTDFILL2_1984 VDD VSS sg13g2_FILL8
XSTDFILL2_1992 VDD VSS sg13g2_FILL8
XSTDFILL2_2000 VDD VSS sg13g2_FILL8
XSTDFILL2_2008 VDD VSS sg13g2_FILL8
XSTDFILL2_2016 VDD VSS sg13g2_FILL8
XSTDFILL2_2024 VDD VSS sg13g2_FILL8
XSTDFILL2_2032 VDD VSS sg13g2_FILL8
XSTDFILL2_2040 VDD VSS sg13g2_FILL8
XSTDFILL2_2048 VDD VSS sg13g2_FILL8
XSTDFILL2_2056 VDD VSS sg13g2_FILL8
XSTDFILL2_2064 VDD VSS sg13g2_FILL8
XSTDFILL2_2072 VDD VSS sg13g2_FILL8
XSTDFILL2_2080 VDD VSS sg13g2_FILL8
XSTDFILL2_2088 VDD VSS sg13g2_FILL8
XSTDFILL2_2096 VDD VSS sg13g2_FILL8
XSTDFILL2_2104 VDD VSS sg13g2_FILL8
XSTDFILL2_2112 VDD VSS sg13g2_FILL8
XSTDFILL2_2120 VDD VSS sg13g2_FILL8
XSTDFILL2_2128 VDD VSS sg13g2_FILL8
XSTDFILL2_2136 VDD VSS sg13g2_FILL8
XSTDFILL2_2144 VDD VSS sg13g2_FILL8
XSTDFILL2_2152 VDD VSS sg13g2_FILL8
XSTDFILL2_2160 VDD VSS sg13g2_FILL8
XSTDFILL2_2168 VDD VSS sg13g2_FILL4
XSTDFILL3_0 VDD VSS sg13g2_FILL8
XSTDFILL3_8 VDD VSS sg13g2_FILL8
XSTDFILL3_16 VDD VSS sg13g2_FILL8
XSTDFILL3_24 VDD VSS sg13g2_FILL8
XSTDFILL3_32 VDD VSS sg13g2_FILL8
XSTDFILL3_40 VDD VSS sg13g2_FILL8
XSTDFILL3_48 VDD VSS sg13g2_FILL8
XSTDFILL3_56 VDD VSS sg13g2_FILL8
XSTDFILL3_64 VDD VSS sg13g2_FILL8
XSTDFILL3_72 VDD VSS sg13g2_FILL8
XSTDFILL3_80 VDD VSS sg13g2_FILL8
XSTDFILL3_88 VDD VSS sg13g2_FILL8
XSTDFILL3_96 VDD VSS sg13g2_FILL8
XSTDFILL3_104 VDD VSS sg13g2_FILL1
XSTDFILL3_1880 VDD VSS sg13g2_FILL8
XSTDFILL3_1888 VDD VSS sg13g2_FILL8
XSTDFILL3_1896 VDD VSS sg13g2_FILL8
XSTDFILL3_1904 VDD VSS sg13g2_FILL8
XSTDFILL3_1912 VDD VSS sg13g2_FILL8
XSTDFILL3_1920 VDD VSS sg13g2_FILL8
XSTDFILL3_1928 VDD VSS sg13g2_FILL8
XSTDFILL3_1936 VDD VSS sg13g2_FILL8
XSTDFILL3_1944 VDD VSS sg13g2_FILL8
XSTDFILL3_1952 VDD VSS sg13g2_FILL8
XSTDFILL3_1960 VDD VSS sg13g2_FILL8
XSTDFILL3_1968 VDD VSS sg13g2_FILL8
XSTDFILL3_1976 VDD VSS sg13g2_FILL8
XSTDFILL3_1984 VDD VSS sg13g2_FILL8
XSTDFILL3_1992 VDD VSS sg13g2_FILL8
XSTDFILL3_2000 VDD VSS sg13g2_FILL8
XSTDFILL3_2008 VDD VSS sg13g2_FILL8
XSTDFILL3_2016 VDD VSS sg13g2_FILL8
XSTDFILL3_2024 VDD VSS sg13g2_FILL8
XSTDFILL3_2032 VDD VSS sg13g2_FILL8
XSTDFILL3_2040 VDD VSS sg13g2_FILL8
XSTDFILL3_2048 VDD VSS sg13g2_FILL8
XSTDFILL3_2056 VDD VSS sg13g2_FILL8
XSTDFILL3_2064 VDD VSS sg13g2_FILL8
XSTDFILL3_2072 VDD VSS sg13g2_FILL8
XSTDFILL3_2080 VDD VSS sg13g2_FILL8
XSTDFILL3_2088 VDD VSS sg13g2_FILL8
XSTDFILL3_2096 VDD VSS sg13g2_FILL8
XSTDFILL3_2104 VDD VSS sg13g2_FILL8
XSTDFILL3_2112 VDD VSS sg13g2_FILL8
XSTDFILL3_2120 VDD VSS sg13g2_FILL8
XSTDFILL3_2128 VDD VSS sg13g2_FILL8
XSTDFILL3_2136 VDD VSS sg13g2_FILL8
XSTDFILL3_2144 VDD VSS sg13g2_FILL8
XSTDFILL3_2152 VDD VSS sg13g2_FILL8
XSTDFILL3_2160 VDD VSS sg13g2_FILL8
XSTDFILL3_2168 VDD VSS sg13g2_FILL4
XSTDFILL4_0 VDD VSS sg13g2_FILL8
XSTDFILL4_8 VDD VSS sg13g2_FILL8
XSTDFILL4_16 VDD VSS sg13g2_FILL8
XSTDFILL4_24 VDD VSS sg13g2_FILL8
XSTDFILL4_32 VDD VSS sg13g2_FILL8
XSTDFILL4_40 VDD VSS sg13g2_FILL8
XSTDFILL4_48 VDD VSS sg13g2_FILL8
XSTDFILL4_56 VDD VSS sg13g2_FILL8
XSTDFILL4_64 VDD VSS sg13g2_FILL8
XSTDFILL4_72 VDD VSS sg13g2_FILL8
XSTDFILL4_80 VDD VSS sg13g2_FILL8
XSTDFILL4_88 VDD VSS sg13g2_FILL8
XSTDFILL4_96 VDD VSS sg13g2_FILL8
XSTDFILL4_104 VDD VSS sg13g2_FILL1
XSTDFILL4_1880 VDD VSS sg13g2_FILL8
XSTDFILL4_1888 VDD VSS sg13g2_FILL8
XSTDFILL4_1896 VDD VSS sg13g2_FILL8
XSTDFILL4_1904 VDD VSS sg13g2_FILL8
XSTDFILL4_1912 VDD VSS sg13g2_FILL8
XSTDFILL4_1920 VDD VSS sg13g2_FILL8
XSTDFILL4_1928 VDD VSS sg13g2_FILL8
XSTDFILL4_1936 VDD VSS sg13g2_FILL8
XSTDFILL4_1944 VDD VSS sg13g2_FILL8
XSTDFILL4_1952 VDD VSS sg13g2_FILL8
XSTDFILL4_1960 VDD VSS sg13g2_FILL8
XSTDFILL4_1968 VDD VSS sg13g2_FILL8
XSTDFILL4_1976 VDD VSS sg13g2_FILL8
XSTDFILL4_1984 VDD VSS sg13g2_FILL8
XSTDFILL4_1992 VDD VSS sg13g2_FILL8
XSTDFILL4_2000 VDD VSS sg13g2_FILL8
XSTDFILL4_2008 VDD VSS sg13g2_FILL8
XSTDFILL4_2016 VDD VSS sg13g2_FILL8
XSTDFILL4_2024 VDD VSS sg13g2_FILL8
XSTDFILL4_2032 VDD VSS sg13g2_FILL8
XSTDFILL4_2040 VDD VSS sg13g2_FILL8
XSTDFILL4_2048 VDD VSS sg13g2_FILL8
XSTDFILL4_2056 VDD VSS sg13g2_FILL8
XSTDFILL4_2064 VDD VSS sg13g2_FILL8
XSTDFILL4_2072 VDD VSS sg13g2_FILL8
XSTDFILL4_2080 VDD VSS sg13g2_FILL8
XSTDFILL4_2088 VDD VSS sg13g2_FILL8
XSTDFILL4_2096 VDD VSS sg13g2_FILL8
XSTDFILL4_2104 VDD VSS sg13g2_FILL8
XSTDFILL4_2112 VDD VSS sg13g2_FILL8
XSTDFILL4_2120 VDD VSS sg13g2_FILL8
XSTDFILL4_2128 VDD VSS sg13g2_FILL8
XSTDFILL4_2136 VDD VSS sg13g2_FILL8
XSTDFILL4_2144 VDD VSS sg13g2_FILL8
XSTDFILL4_2152 VDD VSS sg13g2_FILL8
XSTDFILL4_2160 VDD VSS sg13g2_FILL8
XSTDFILL4_2168 VDD VSS sg13g2_FILL4
XSTDFILL5_0 VDD VSS sg13g2_FILL8
XSTDFILL5_8 VDD VSS sg13g2_FILL8
XSTDFILL5_16 VDD VSS sg13g2_FILL8
XSTDFILL5_24 VDD VSS sg13g2_FILL8
XSTDFILL5_32 VDD VSS sg13g2_FILL8
XSTDFILL5_40 VDD VSS sg13g2_FILL8
XSTDFILL5_48 VDD VSS sg13g2_FILL8
XSTDFILL5_56 VDD VSS sg13g2_FILL8
XSTDFILL5_64 VDD VSS sg13g2_FILL8
XSTDFILL5_72 VDD VSS sg13g2_FILL8
XSTDFILL5_80 VDD VSS sg13g2_FILL8
XSTDFILL5_88 VDD VSS sg13g2_FILL8
XSTDFILL5_96 VDD VSS sg13g2_FILL8
XSTDFILL5_104 VDD VSS sg13g2_FILL1
XSTDFILL5_1880 VDD VSS sg13g2_FILL8
XSTDFILL5_1888 VDD VSS sg13g2_FILL8
XSTDFILL5_1896 VDD VSS sg13g2_FILL8
XSTDFILL5_1904 VDD VSS sg13g2_FILL8
XSTDFILL5_1912 VDD VSS sg13g2_FILL8
XSTDFILL5_1920 VDD VSS sg13g2_FILL8
XSTDFILL5_1928 VDD VSS sg13g2_FILL8
XSTDFILL5_1936 VDD VSS sg13g2_FILL8
XSTDFILL5_1944 VDD VSS sg13g2_FILL8
XSTDFILL5_1952 VDD VSS sg13g2_FILL8
XSTDFILL5_1960 VDD VSS sg13g2_FILL8
XSTDFILL5_1968 VDD VSS sg13g2_FILL8
XSTDFILL5_1976 VDD VSS sg13g2_FILL8
XSTDFILL5_1984 VDD VSS sg13g2_FILL8
XSTDFILL5_1992 VDD VSS sg13g2_FILL8
XSTDFILL5_2000 VDD VSS sg13g2_FILL8
XSTDFILL5_2008 VDD VSS sg13g2_FILL8
XSTDFILL5_2016 VDD VSS sg13g2_FILL8
XSTDFILL5_2024 VDD VSS sg13g2_FILL8
XSTDFILL5_2032 VDD VSS sg13g2_FILL8
XSTDFILL5_2040 VDD VSS sg13g2_FILL8
XSTDFILL5_2048 VDD VSS sg13g2_FILL8
XSTDFILL5_2056 VDD VSS sg13g2_FILL8
XSTDFILL5_2064 VDD VSS sg13g2_FILL8
XSTDFILL5_2072 VDD VSS sg13g2_FILL8
XSTDFILL5_2080 VDD VSS sg13g2_FILL8
XSTDFILL5_2088 VDD VSS sg13g2_FILL8
XSTDFILL5_2096 VDD VSS sg13g2_FILL8
XSTDFILL5_2104 VDD VSS sg13g2_FILL8
XSTDFILL5_2112 VDD VSS sg13g2_FILL8
XSTDFILL5_2120 VDD VSS sg13g2_FILL8
XSTDFILL5_2128 VDD VSS sg13g2_FILL8
XSTDFILL5_2136 VDD VSS sg13g2_FILL8
XSTDFILL5_2144 VDD VSS sg13g2_FILL8
XSTDFILL5_2152 VDD VSS sg13g2_FILL8
XSTDFILL5_2160 VDD VSS sg13g2_FILL8
XSTDFILL5_2168 VDD VSS sg13g2_FILL4
XSTDFILL6_0 VDD VSS sg13g2_FILL8
XSTDFILL6_8 VDD VSS sg13g2_FILL8
XSTDFILL6_16 VDD VSS sg13g2_FILL8
XSTDFILL6_24 VDD VSS sg13g2_FILL8
XSTDFILL6_32 VDD VSS sg13g2_FILL8
XSTDFILL6_40 VDD VSS sg13g2_FILL8
XSTDFILL6_48 VDD VSS sg13g2_FILL8
XSTDFILL6_56 VDD VSS sg13g2_FILL8
XSTDFILL6_64 VDD VSS sg13g2_FILL8
XSTDFILL6_72 VDD VSS sg13g2_FILL8
XSTDFILL6_80 VDD VSS sg13g2_FILL8
XSTDFILL6_88 VDD VSS sg13g2_FILL8
XSTDFILL6_96 VDD VSS sg13g2_FILL8
XSTDFILL6_104 VDD VSS sg13g2_FILL1
XSTDFILL6_1880 VDD VSS sg13g2_FILL8
XSTDFILL6_1888 VDD VSS sg13g2_FILL8
XSTDFILL6_1896 VDD VSS sg13g2_FILL8
XSTDFILL6_1904 VDD VSS sg13g2_FILL8
XSTDFILL6_1912 VDD VSS sg13g2_FILL8
XSTDFILL6_1920 VDD VSS sg13g2_FILL8
XSTDFILL6_1928 VDD VSS sg13g2_FILL8
XSTDFILL6_1936 VDD VSS sg13g2_FILL8
XSTDFILL6_1944 VDD VSS sg13g2_FILL8
XSTDFILL6_1952 VDD VSS sg13g2_FILL8
XSTDFILL6_1960 VDD VSS sg13g2_FILL8
XSTDFILL6_1968 VDD VSS sg13g2_FILL8
XSTDFILL6_1976 VDD VSS sg13g2_FILL8
XSTDFILL6_1984 VDD VSS sg13g2_FILL8
XSTDFILL6_1992 VDD VSS sg13g2_FILL8
XSTDFILL6_2000 VDD VSS sg13g2_FILL8
XSTDFILL6_2008 VDD VSS sg13g2_FILL8
XSTDFILL6_2016 VDD VSS sg13g2_FILL8
XSTDFILL6_2024 VDD VSS sg13g2_FILL8
XSTDFILL6_2032 VDD VSS sg13g2_FILL8
XSTDFILL6_2040 VDD VSS sg13g2_FILL8
XSTDFILL6_2048 VDD VSS sg13g2_FILL8
XSTDFILL6_2056 VDD VSS sg13g2_FILL8
XSTDFILL6_2064 VDD VSS sg13g2_FILL8
XSTDFILL6_2072 VDD VSS sg13g2_FILL8
XSTDFILL6_2080 VDD VSS sg13g2_FILL8
XSTDFILL6_2088 VDD VSS sg13g2_FILL8
XSTDFILL6_2096 VDD VSS sg13g2_FILL8
XSTDFILL6_2104 VDD VSS sg13g2_FILL8
XSTDFILL6_2112 VDD VSS sg13g2_FILL8
XSTDFILL6_2120 VDD VSS sg13g2_FILL8
XSTDFILL6_2128 VDD VSS sg13g2_FILL8
XSTDFILL6_2136 VDD VSS sg13g2_FILL8
XSTDFILL6_2144 VDD VSS sg13g2_FILL8
XSTDFILL6_2152 VDD VSS sg13g2_FILL8
XSTDFILL6_2160 VDD VSS sg13g2_FILL8
XSTDFILL6_2168 VDD VSS sg13g2_FILL4
XSTDFILL7_0 VDD VSS sg13g2_FILL8
XSTDFILL7_8 VDD VSS sg13g2_FILL8
XSTDFILL7_16 VDD VSS sg13g2_FILL8
XSTDFILL7_24 VDD VSS sg13g2_FILL8
XSTDFILL7_32 VDD VSS sg13g2_FILL8
XSTDFILL7_40 VDD VSS sg13g2_FILL8
XSTDFILL7_48 VDD VSS sg13g2_FILL8
XSTDFILL7_56 VDD VSS sg13g2_FILL8
XSTDFILL7_64 VDD VSS sg13g2_FILL8
XSTDFILL7_72 VDD VSS sg13g2_FILL8
XSTDFILL7_80 VDD VSS sg13g2_FILL8
XSTDFILL7_88 VDD VSS sg13g2_FILL8
XSTDFILL7_96 VDD VSS sg13g2_FILL8
XSTDFILL7_104 VDD VSS sg13g2_FILL1
XSTDFILL7_1880 VDD VSS sg13g2_FILL8
XSTDFILL7_1888 VDD VSS sg13g2_FILL8
XSTDFILL7_1896 VDD VSS sg13g2_FILL8
XSTDFILL7_1904 VDD VSS sg13g2_FILL8
XSTDFILL7_1912 VDD VSS sg13g2_FILL8
XSTDFILL7_1920 VDD VSS sg13g2_FILL8
XSTDFILL7_1928 VDD VSS sg13g2_FILL8
XSTDFILL7_1936 VDD VSS sg13g2_FILL8
XSTDFILL7_1944 VDD VSS sg13g2_FILL8
XSTDFILL7_1952 VDD VSS sg13g2_FILL8
XSTDFILL7_1960 VDD VSS sg13g2_FILL8
XSTDFILL7_1968 VDD VSS sg13g2_FILL8
XSTDFILL7_1976 VDD VSS sg13g2_FILL8
XSTDFILL7_1984 VDD VSS sg13g2_FILL8
XSTDFILL7_1992 VDD VSS sg13g2_FILL8
XSTDFILL7_2000 VDD VSS sg13g2_FILL8
XSTDFILL7_2008 VDD VSS sg13g2_FILL8
XSTDFILL7_2016 VDD VSS sg13g2_FILL8
XSTDFILL7_2024 VDD VSS sg13g2_FILL8
XSTDFILL7_2032 VDD VSS sg13g2_FILL8
XSTDFILL7_2040 VDD VSS sg13g2_FILL8
XSTDFILL7_2048 VDD VSS sg13g2_FILL8
XSTDFILL7_2056 VDD VSS sg13g2_FILL8
XSTDFILL7_2064 VDD VSS sg13g2_FILL8
XSTDFILL7_2072 VDD VSS sg13g2_FILL8
XSTDFILL7_2080 VDD VSS sg13g2_FILL8
XSTDFILL7_2088 VDD VSS sg13g2_FILL8
XSTDFILL7_2096 VDD VSS sg13g2_FILL8
XSTDFILL7_2104 VDD VSS sg13g2_FILL8
XSTDFILL7_2112 VDD VSS sg13g2_FILL8
XSTDFILL7_2120 VDD VSS sg13g2_FILL8
XSTDFILL7_2128 VDD VSS sg13g2_FILL8
XSTDFILL7_2136 VDD VSS sg13g2_FILL8
XSTDFILL7_2144 VDD VSS sg13g2_FILL8
XSTDFILL7_2152 VDD VSS sg13g2_FILL8
XSTDFILL7_2160 VDD VSS sg13g2_FILL8
XSTDFILL7_2168 VDD VSS sg13g2_FILL4
XSTDFILL8_0 VDD VSS sg13g2_FILL8
XSTDFILL8_8 VDD VSS sg13g2_FILL8
XSTDFILL8_16 VDD VSS sg13g2_FILL8
XSTDFILL8_24 VDD VSS sg13g2_FILL8
XSTDFILL8_32 VDD VSS sg13g2_FILL8
XSTDFILL8_40 VDD VSS sg13g2_FILL8
XSTDFILL8_48 VDD VSS sg13g2_FILL8
XSTDFILL8_56 VDD VSS sg13g2_FILL8
XSTDFILL8_64 VDD VSS sg13g2_FILL8
XSTDFILL8_72 VDD VSS sg13g2_FILL8
XSTDFILL8_80 VDD VSS sg13g2_FILL8
XSTDFILL8_88 VDD VSS sg13g2_FILL8
XSTDFILL8_96 VDD VSS sg13g2_FILL8
XSTDFILL8_104 VDD VSS sg13g2_FILL1
XSTDFILL8_1880 VDD VSS sg13g2_FILL8
XSTDFILL8_1888 VDD VSS sg13g2_FILL8
XSTDFILL8_1896 VDD VSS sg13g2_FILL8
XSTDFILL8_1904 VDD VSS sg13g2_FILL8
XSTDFILL8_1912 VDD VSS sg13g2_FILL8
XSTDFILL8_1920 VDD VSS sg13g2_FILL8
XSTDFILL8_1928 VDD VSS sg13g2_FILL8
XSTDFILL8_1936 VDD VSS sg13g2_FILL8
XSTDFILL8_1944 VDD VSS sg13g2_FILL8
XSTDFILL8_1952 VDD VSS sg13g2_FILL8
XSTDFILL8_1960 VDD VSS sg13g2_FILL8
XSTDFILL8_1968 VDD VSS sg13g2_FILL8
XSTDFILL8_1976 VDD VSS sg13g2_FILL8
XSTDFILL8_1984 VDD VSS sg13g2_FILL8
XSTDFILL8_1992 VDD VSS sg13g2_FILL8
XSTDFILL8_2000 VDD VSS sg13g2_FILL8
XSTDFILL8_2008 VDD VSS sg13g2_FILL8
XSTDFILL8_2016 VDD VSS sg13g2_FILL8
XSTDFILL8_2024 VDD VSS sg13g2_FILL8
XSTDFILL8_2032 VDD VSS sg13g2_FILL8
XSTDFILL8_2040 VDD VSS sg13g2_FILL8
XSTDFILL8_2048 VDD VSS sg13g2_FILL8
XSTDFILL8_2056 VDD VSS sg13g2_FILL8
XSTDFILL8_2064 VDD VSS sg13g2_FILL8
XSTDFILL8_2072 VDD VSS sg13g2_FILL8
XSTDFILL8_2080 VDD VSS sg13g2_FILL8
XSTDFILL8_2088 VDD VSS sg13g2_FILL8
XSTDFILL8_2096 VDD VSS sg13g2_FILL8
XSTDFILL8_2104 VDD VSS sg13g2_FILL8
XSTDFILL8_2112 VDD VSS sg13g2_FILL8
XSTDFILL8_2120 VDD VSS sg13g2_FILL8
XSTDFILL8_2128 VDD VSS sg13g2_FILL8
XSTDFILL8_2136 VDD VSS sg13g2_FILL8
XSTDFILL8_2144 VDD VSS sg13g2_FILL8
XSTDFILL8_2152 VDD VSS sg13g2_FILL8
XSTDFILL8_2160 VDD VSS sg13g2_FILL8
XSTDFILL8_2168 VDD VSS sg13g2_FILL4
XSTDFILL9_0 VDD VSS sg13g2_FILL8
XSTDFILL9_8 VDD VSS sg13g2_FILL8
XSTDFILL9_16 VDD VSS sg13g2_FILL8
XSTDFILL9_24 VDD VSS sg13g2_FILL8
XSTDFILL9_32 VDD VSS sg13g2_FILL8
XSTDFILL9_40 VDD VSS sg13g2_FILL8
XSTDFILL9_48 VDD VSS sg13g2_FILL8
XSTDFILL9_56 VDD VSS sg13g2_FILL8
XSTDFILL9_64 VDD VSS sg13g2_FILL8
XSTDFILL9_72 VDD VSS sg13g2_FILL8
XSTDFILL9_80 VDD VSS sg13g2_FILL8
XSTDFILL9_88 VDD VSS sg13g2_FILL8
XSTDFILL9_96 VDD VSS sg13g2_FILL8
XSTDFILL9_104 VDD VSS sg13g2_FILL1
XSTDFILL9_1880 VDD VSS sg13g2_FILL8
XSTDFILL9_1888 VDD VSS sg13g2_FILL8
XSTDFILL9_1896 VDD VSS sg13g2_FILL8
XSTDFILL9_1904 VDD VSS sg13g2_FILL8
XSTDFILL9_1912 VDD VSS sg13g2_FILL8
XSTDFILL9_1920 VDD VSS sg13g2_FILL8
XSTDFILL9_1928 VDD VSS sg13g2_FILL8
XSTDFILL9_1936 VDD VSS sg13g2_FILL8
XSTDFILL9_1944 VDD VSS sg13g2_FILL8
XSTDFILL9_1952 VDD VSS sg13g2_FILL8
XSTDFILL9_1960 VDD VSS sg13g2_FILL8
XSTDFILL9_1968 VDD VSS sg13g2_FILL8
XSTDFILL9_1976 VDD VSS sg13g2_FILL8
XSTDFILL9_1984 VDD VSS sg13g2_FILL8
XSTDFILL9_1992 VDD VSS sg13g2_FILL8
XSTDFILL9_2000 VDD VSS sg13g2_FILL8
XSTDFILL9_2008 VDD VSS sg13g2_FILL8
XSTDFILL9_2016 VDD VSS sg13g2_FILL8
XSTDFILL9_2024 VDD VSS sg13g2_FILL8
XSTDFILL9_2032 VDD VSS sg13g2_FILL8
XSTDFILL9_2040 VDD VSS sg13g2_FILL8
XSTDFILL9_2048 VDD VSS sg13g2_FILL8
XSTDFILL9_2056 VDD VSS sg13g2_FILL8
XSTDFILL9_2064 VDD VSS sg13g2_FILL8
XSTDFILL9_2072 VDD VSS sg13g2_FILL8
XSTDFILL9_2080 VDD VSS sg13g2_FILL8
XSTDFILL9_2088 VDD VSS sg13g2_FILL8
XSTDFILL9_2096 VDD VSS sg13g2_FILL8
XSTDFILL9_2104 VDD VSS sg13g2_FILL8
XSTDFILL9_2112 VDD VSS sg13g2_FILL8
XSTDFILL9_2120 VDD VSS sg13g2_FILL8
XSTDFILL9_2128 VDD VSS sg13g2_FILL8
XSTDFILL9_2136 VDD VSS sg13g2_FILL8
XSTDFILL9_2144 VDD VSS sg13g2_FILL8
XSTDFILL9_2152 VDD VSS sg13g2_FILL8
XSTDFILL9_2160 VDD VSS sg13g2_FILL8
XSTDFILL9_2168 VDD VSS sg13g2_FILL4
XSTDFILL10_0 VDD VSS sg13g2_FILL8
XSTDFILL10_8 VDD VSS sg13g2_FILL8
XSTDFILL10_16 VDD VSS sg13g2_FILL8
XSTDFILL10_24 VDD VSS sg13g2_FILL8
XSTDFILL10_32 VDD VSS sg13g2_FILL8
XSTDFILL10_40 VDD VSS sg13g2_FILL8
XSTDFILL10_48 VDD VSS sg13g2_FILL8
XSTDFILL10_56 VDD VSS sg13g2_FILL8
XSTDFILL10_64 VDD VSS sg13g2_FILL8
XSTDFILL10_72 VDD VSS sg13g2_FILL8
XSTDFILL10_80 VDD VSS sg13g2_FILL8
XSTDFILL10_88 VDD VSS sg13g2_FILL8
XSTDFILL10_96 VDD VSS sg13g2_FILL8
XSTDFILL10_104 VDD VSS sg13g2_FILL1
XSTDFILL10_1880 VDD VSS sg13g2_FILL8
XSTDFILL10_1888 VDD VSS sg13g2_FILL8
XSTDFILL10_1896 VDD VSS sg13g2_FILL8
XSTDFILL10_1904 VDD VSS sg13g2_FILL8
XSTDFILL10_1912 VDD VSS sg13g2_FILL8
XSTDFILL10_1920 VDD VSS sg13g2_FILL8
XSTDFILL10_1928 VDD VSS sg13g2_FILL8
XSTDFILL10_1936 VDD VSS sg13g2_FILL8
XSTDFILL10_1944 VDD VSS sg13g2_FILL8
XSTDFILL10_1952 VDD VSS sg13g2_FILL8
XSTDFILL10_1960 VDD VSS sg13g2_FILL8
XSTDFILL10_1968 VDD VSS sg13g2_FILL8
XSTDFILL10_1976 VDD VSS sg13g2_FILL8
XSTDFILL10_1984 VDD VSS sg13g2_FILL8
XSTDFILL10_1992 VDD VSS sg13g2_FILL8
XSTDFILL10_2000 VDD VSS sg13g2_FILL8
XSTDFILL10_2008 VDD VSS sg13g2_FILL8
XSTDFILL10_2016 VDD VSS sg13g2_FILL8
XSTDFILL10_2024 VDD VSS sg13g2_FILL8
XSTDFILL10_2032 VDD VSS sg13g2_FILL8
XSTDFILL10_2040 VDD VSS sg13g2_FILL8
XSTDFILL10_2048 VDD VSS sg13g2_FILL8
XSTDFILL10_2056 VDD VSS sg13g2_FILL8
XSTDFILL10_2064 VDD VSS sg13g2_FILL8
XSTDFILL10_2072 VDD VSS sg13g2_FILL8
XSTDFILL10_2080 VDD VSS sg13g2_FILL8
XSTDFILL10_2088 VDD VSS sg13g2_FILL8
XSTDFILL10_2096 VDD VSS sg13g2_FILL8
XSTDFILL10_2104 VDD VSS sg13g2_FILL8
XSTDFILL10_2112 VDD VSS sg13g2_FILL8
XSTDFILL10_2120 VDD VSS sg13g2_FILL8
XSTDFILL10_2128 VDD VSS sg13g2_FILL8
XSTDFILL10_2136 VDD VSS sg13g2_FILL8
XSTDFILL10_2144 VDD VSS sg13g2_FILL8
XSTDFILL10_2152 VDD VSS sg13g2_FILL8
XSTDFILL10_2160 VDD VSS sg13g2_FILL8
XSTDFILL10_2168 VDD VSS sg13g2_FILL4
XSTDFILL11_0 VDD VSS sg13g2_FILL8
XSTDFILL11_8 VDD VSS sg13g2_FILL8
XSTDFILL11_16 VDD VSS sg13g2_FILL8
XSTDFILL11_24 VDD VSS sg13g2_FILL8
XSTDFILL11_32 VDD VSS sg13g2_FILL8
XSTDFILL11_40 VDD VSS sg13g2_FILL8
XSTDFILL11_48 VDD VSS sg13g2_FILL8
XSTDFILL11_56 VDD VSS sg13g2_FILL8
XSTDFILL11_64 VDD VSS sg13g2_FILL8
XSTDFILL11_72 VDD VSS sg13g2_FILL8
XSTDFILL11_80 VDD VSS sg13g2_FILL8
XSTDFILL11_88 VDD VSS sg13g2_FILL8
XSTDFILL11_96 VDD VSS sg13g2_FILL8
XSTDFILL11_104 VDD VSS sg13g2_FILL1
XSTDFILL11_1880 VDD VSS sg13g2_FILL8
XSTDFILL11_1888 VDD VSS sg13g2_FILL8
XSTDFILL11_1896 VDD VSS sg13g2_FILL8
XSTDFILL11_1904 VDD VSS sg13g2_FILL8
XSTDFILL11_1912 VDD VSS sg13g2_FILL8
XSTDFILL11_1920 VDD VSS sg13g2_FILL8
XSTDFILL11_1928 VDD VSS sg13g2_FILL8
XSTDFILL11_1936 VDD VSS sg13g2_FILL8
XSTDFILL11_1944 VDD VSS sg13g2_FILL8
XSTDFILL11_1952 VDD VSS sg13g2_FILL8
XSTDFILL11_1960 VDD VSS sg13g2_FILL8
XSTDFILL11_1968 VDD VSS sg13g2_FILL8
XSTDFILL11_1976 VDD VSS sg13g2_FILL8
XSTDFILL11_1984 VDD VSS sg13g2_FILL8
XSTDFILL11_1992 VDD VSS sg13g2_FILL8
XSTDFILL11_2000 VDD VSS sg13g2_FILL8
XSTDFILL11_2008 VDD VSS sg13g2_FILL8
XSTDFILL11_2016 VDD VSS sg13g2_FILL8
XSTDFILL11_2024 VDD VSS sg13g2_FILL8
XSTDFILL11_2032 VDD VSS sg13g2_FILL8
XSTDFILL11_2040 VDD VSS sg13g2_FILL8
XSTDFILL11_2048 VDD VSS sg13g2_FILL8
XSTDFILL11_2056 VDD VSS sg13g2_FILL8
XSTDFILL11_2064 VDD VSS sg13g2_FILL8
XSTDFILL11_2072 VDD VSS sg13g2_FILL8
XSTDFILL11_2080 VDD VSS sg13g2_FILL8
XSTDFILL11_2088 VDD VSS sg13g2_FILL8
XSTDFILL11_2096 VDD VSS sg13g2_FILL8
XSTDFILL11_2104 VDD VSS sg13g2_FILL8
XSTDFILL11_2112 VDD VSS sg13g2_FILL8
XSTDFILL11_2120 VDD VSS sg13g2_FILL8
XSTDFILL11_2128 VDD VSS sg13g2_FILL8
XSTDFILL11_2136 VDD VSS sg13g2_FILL8
XSTDFILL11_2144 VDD VSS sg13g2_FILL8
XSTDFILL11_2152 VDD VSS sg13g2_FILL8
XSTDFILL11_2160 VDD VSS sg13g2_FILL8
XSTDFILL11_2168 VDD VSS sg13g2_FILL4
XSTDFILL12_0 VDD VSS sg13g2_FILL8
XSTDFILL12_8 VDD VSS sg13g2_FILL8
XSTDFILL12_16 VDD VSS sg13g2_FILL8
XSTDFILL12_24 VDD VSS sg13g2_FILL8
XSTDFILL12_32 VDD VSS sg13g2_FILL8
XSTDFILL12_40 VDD VSS sg13g2_FILL8
XSTDFILL12_48 VDD VSS sg13g2_FILL8
XSTDFILL12_56 VDD VSS sg13g2_FILL8
XSTDFILL12_64 VDD VSS sg13g2_FILL8
XSTDFILL12_72 VDD VSS sg13g2_FILL8
XSTDFILL12_80 VDD VSS sg13g2_FILL8
XSTDFILL12_88 VDD VSS sg13g2_FILL8
XSTDFILL12_96 VDD VSS sg13g2_FILL8
XSTDFILL12_104 VDD VSS sg13g2_FILL1
XSTDFILL12_1880 VDD VSS sg13g2_FILL8
XSTDFILL12_1888 VDD VSS sg13g2_FILL8
XSTDFILL12_1896 VDD VSS sg13g2_FILL8
XSTDFILL12_1904 VDD VSS sg13g2_FILL8
XSTDFILL12_1912 VDD VSS sg13g2_FILL8
XSTDFILL12_1920 VDD VSS sg13g2_FILL8
XSTDFILL12_1928 VDD VSS sg13g2_FILL8
XSTDFILL12_1936 VDD VSS sg13g2_FILL8
XSTDFILL12_1944 VDD VSS sg13g2_FILL8
XSTDFILL12_1952 VDD VSS sg13g2_FILL8
XSTDFILL12_1960 VDD VSS sg13g2_FILL8
XSTDFILL12_1968 VDD VSS sg13g2_FILL8
XSTDFILL12_1976 VDD VSS sg13g2_FILL8
XSTDFILL12_1984 VDD VSS sg13g2_FILL8
XSTDFILL12_1992 VDD VSS sg13g2_FILL8
XSTDFILL12_2000 VDD VSS sg13g2_FILL8
XSTDFILL12_2008 VDD VSS sg13g2_FILL8
XSTDFILL12_2016 VDD VSS sg13g2_FILL8
XSTDFILL12_2024 VDD VSS sg13g2_FILL8
XSTDFILL12_2032 VDD VSS sg13g2_FILL8
XSTDFILL12_2040 VDD VSS sg13g2_FILL8
XSTDFILL12_2048 VDD VSS sg13g2_FILL8
XSTDFILL12_2056 VDD VSS sg13g2_FILL8
XSTDFILL12_2064 VDD VSS sg13g2_FILL8
XSTDFILL12_2072 VDD VSS sg13g2_FILL8
XSTDFILL12_2080 VDD VSS sg13g2_FILL8
XSTDFILL12_2088 VDD VSS sg13g2_FILL8
XSTDFILL12_2096 VDD VSS sg13g2_FILL8
XSTDFILL12_2104 VDD VSS sg13g2_FILL8
XSTDFILL12_2112 VDD VSS sg13g2_FILL8
XSTDFILL12_2120 VDD VSS sg13g2_FILL8
XSTDFILL12_2128 VDD VSS sg13g2_FILL8
XSTDFILL12_2136 VDD VSS sg13g2_FILL8
XSTDFILL12_2144 VDD VSS sg13g2_FILL8
XSTDFILL12_2152 VDD VSS sg13g2_FILL8
XSTDFILL12_2160 VDD VSS sg13g2_FILL8
XSTDFILL12_2168 VDD VSS sg13g2_FILL4
XSTDFILL13_0 VDD VSS sg13g2_FILL8
XSTDFILL13_8 VDD VSS sg13g2_FILL8
XSTDFILL13_16 VDD VSS sg13g2_FILL8
XSTDFILL13_24 VDD VSS sg13g2_FILL8
XSTDFILL13_32 VDD VSS sg13g2_FILL8
XSTDFILL13_40 VDD VSS sg13g2_FILL8
XSTDFILL13_48 VDD VSS sg13g2_FILL8
XSTDFILL13_56 VDD VSS sg13g2_FILL8
XSTDFILL13_64 VDD VSS sg13g2_FILL8
XSTDFILL13_72 VDD VSS sg13g2_FILL8
XSTDFILL13_80 VDD VSS sg13g2_FILL8
XSTDFILL13_88 VDD VSS sg13g2_FILL8
XSTDFILL13_96 VDD VSS sg13g2_FILL8
XSTDFILL13_104 VDD VSS sg13g2_FILL1
XSTDFILL13_1880 VDD VSS sg13g2_FILL8
XSTDFILL13_1888 VDD VSS sg13g2_FILL8
XSTDFILL13_1896 VDD VSS sg13g2_FILL8
XSTDFILL13_1904 VDD VSS sg13g2_FILL8
XSTDFILL13_1912 VDD VSS sg13g2_FILL8
XSTDFILL13_1920 VDD VSS sg13g2_FILL8
XSTDFILL13_1928 VDD VSS sg13g2_FILL8
XSTDFILL13_1936 VDD VSS sg13g2_FILL8
XSTDFILL13_1944 VDD VSS sg13g2_FILL8
XSTDFILL13_1952 VDD VSS sg13g2_FILL8
XSTDFILL13_1960 VDD VSS sg13g2_FILL8
XSTDFILL13_1968 VDD VSS sg13g2_FILL8
XSTDFILL13_1976 VDD VSS sg13g2_FILL8
XSTDFILL13_1984 VDD VSS sg13g2_FILL8
XSTDFILL13_1992 VDD VSS sg13g2_FILL8
XSTDFILL13_2000 VDD VSS sg13g2_FILL8
XSTDFILL13_2008 VDD VSS sg13g2_FILL8
XSTDFILL13_2016 VDD VSS sg13g2_FILL8
XSTDFILL13_2024 VDD VSS sg13g2_FILL8
XSTDFILL13_2032 VDD VSS sg13g2_FILL8
XSTDFILL13_2040 VDD VSS sg13g2_FILL8
XSTDFILL13_2048 VDD VSS sg13g2_FILL8
XSTDFILL13_2056 VDD VSS sg13g2_FILL8
XSTDFILL13_2064 VDD VSS sg13g2_FILL8
XSTDFILL13_2072 VDD VSS sg13g2_FILL8
XSTDFILL13_2080 VDD VSS sg13g2_FILL8
XSTDFILL13_2088 VDD VSS sg13g2_FILL8
XSTDFILL13_2096 VDD VSS sg13g2_FILL8
XSTDFILL13_2104 VDD VSS sg13g2_FILL8
XSTDFILL13_2112 VDD VSS sg13g2_FILL8
XSTDFILL13_2120 VDD VSS sg13g2_FILL8
XSTDFILL13_2128 VDD VSS sg13g2_FILL8
XSTDFILL13_2136 VDD VSS sg13g2_FILL8
XSTDFILL13_2144 VDD VSS sg13g2_FILL8
XSTDFILL13_2152 VDD VSS sg13g2_FILL8
XSTDFILL13_2160 VDD VSS sg13g2_FILL8
XSTDFILL13_2168 VDD VSS sg13g2_FILL4
XSTDFILL14_0 VDD VSS sg13g2_FILL8
XSTDFILL14_8 VDD VSS sg13g2_FILL8
XSTDFILL14_16 VDD VSS sg13g2_FILL8
XSTDFILL14_24 VDD VSS sg13g2_FILL8
XSTDFILL14_32 VDD VSS sg13g2_FILL8
XSTDFILL14_40 VDD VSS sg13g2_FILL8
XSTDFILL14_48 VDD VSS sg13g2_FILL8
XSTDFILL14_56 VDD VSS sg13g2_FILL8
XSTDFILL14_64 VDD VSS sg13g2_FILL8
XSTDFILL14_72 VDD VSS sg13g2_FILL8
XSTDFILL14_80 VDD VSS sg13g2_FILL8
XSTDFILL14_88 VDD VSS sg13g2_FILL8
XSTDFILL14_96 VDD VSS sg13g2_FILL8
XSTDFILL14_104 VDD VSS sg13g2_FILL1
XSTDFILL14_1880 VDD VSS sg13g2_FILL8
XSTDFILL14_1888 VDD VSS sg13g2_FILL8
XSTDFILL14_1896 VDD VSS sg13g2_FILL8
XSTDFILL14_1904 VDD VSS sg13g2_FILL8
XSTDFILL14_1912 VDD VSS sg13g2_FILL8
XSTDFILL14_1920 VDD VSS sg13g2_FILL8
XSTDFILL14_1928 VDD VSS sg13g2_FILL8
XSTDFILL14_1936 VDD VSS sg13g2_FILL8
XSTDFILL14_1944 VDD VSS sg13g2_FILL8
XSTDFILL14_1952 VDD VSS sg13g2_FILL8
XSTDFILL14_1960 VDD VSS sg13g2_FILL8
XSTDFILL14_1968 VDD VSS sg13g2_FILL8
XSTDFILL14_1976 VDD VSS sg13g2_FILL8
XSTDFILL14_1984 VDD VSS sg13g2_FILL8
XSTDFILL14_1992 VDD VSS sg13g2_FILL8
XSTDFILL14_2000 VDD VSS sg13g2_FILL8
XSTDFILL14_2008 VDD VSS sg13g2_FILL8
XSTDFILL14_2016 VDD VSS sg13g2_FILL8
XSTDFILL14_2024 VDD VSS sg13g2_FILL8
XSTDFILL14_2032 VDD VSS sg13g2_FILL8
XSTDFILL14_2040 VDD VSS sg13g2_FILL8
XSTDFILL14_2048 VDD VSS sg13g2_FILL8
XSTDFILL14_2056 VDD VSS sg13g2_FILL8
XSTDFILL14_2064 VDD VSS sg13g2_FILL8
XSTDFILL14_2072 VDD VSS sg13g2_FILL8
XSTDFILL14_2080 VDD VSS sg13g2_FILL8
XSTDFILL14_2088 VDD VSS sg13g2_FILL8
XSTDFILL14_2096 VDD VSS sg13g2_FILL8
XSTDFILL14_2104 VDD VSS sg13g2_FILL8
XSTDFILL14_2112 VDD VSS sg13g2_FILL8
XSTDFILL14_2120 VDD VSS sg13g2_FILL8
XSTDFILL14_2128 VDD VSS sg13g2_FILL8
XSTDFILL14_2136 VDD VSS sg13g2_FILL8
XSTDFILL14_2144 VDD VSS sg13g2_FILL8
XSTDFILL14_2152 VDD VSS sg13g2_FILL8
XSTDFILL14_2160 VDD VSS sg13g2_FILL8
XSTDFILL14_2168 VDD VSS sg13g2_FILL4
XSTDFILL15_0 VDD VSS sg13g2_FILL8
XSTDFILL15_8 VDD VSS sg13g2_FILL8
XSTDFILL15_16 VDD VSS sg13g2_FILL8
XSTDFILL15_24 VDD VSS sg13g2_FILL8
XSTDFILL15_32 VDD VSS sg13g2_FILL8
XSTDFILL15_40 VDD VSS sg13g2_FILL8
XSTDFILL15_48 VDD VSS sg13g2_FILL8
XSTDFILL15_56 VDD VSS sg13g2_FILL8
XSTDFILL15_64 VDD VSS sg13g2_FILL8
XSTDFILL15_72 VDD VSS sg13g2_FILL8
XSTDFILL15_80 VDD VSS sg13g2_FILL8
XSTDFILL15_88 VDD VSS sg13g2_FILL8
XSTDFILL15_96 VDD VSS sg13g2_FILL8
XSTDFILL15_104 VDD VSS sg13g2_FILL1
XSTDFILL15_1880 VDD VSS sg13g2_FILL8
XSTDFILL15_1888 VDD VSS sg13g2_FILL8
XSTDFILL15_1896 VDD VSS sg13g2_FILL8
XSTDFILL15_1904 VDD VSS sg13g2_FILL8
XSTDFILL15_1912 VDD VSS sg13g2_FILL8
XSTDFILL15_1920 VDD VSS sg13g2_FILL8
XSTDFILL15_1928 VDD VSS sg13g2_FILL8
XSTDFILL15_1936 VDD VSS sg13g2_FILL8
XSTDFILL15_1944 VDD VSS sg13g2_FILL8
XSTDFILL15_1952 VDD VSS sg13g2_FILL8
XSTDFILL15_1960 VDD VSS sg13g2_FILL8
XSTDFILL15_1968 VDD VSS sg13g2_FILL8
XSTDFILL15_1976 VDD VSS sg13g2_FILL8
XSTDFILL15_1984 VDD VSS sg13g2_FILL8
XSTDFILL15_1992 VDD VSS sg13g2_FILL8
XSTDFILL15_2000 VDD VSS sg13g2_FILL8
XSTDFILL15_2008 VDD VSS sg13g2_FILL8
XSTDFILL15_2016 VDD VSS sg13g2_FILL8
XSTDFILL15_2024 VDD VSS sg13g2_FILL8
XSTDFILL15_2032 VDD VSS sg13g2_FILL8
XSTDFILL15_2040 VDD VSS sg13g2_FILL8
XSTDFILL15_2048 VDD VSS sg13g2_FILL8
XSTDFILL15_2056 VDD VSS sg13g2_FILL8
XSTDFILL15_2064 VDD VSS sg13g2_FILL8
XSTDFILL15_2072 VDD VSS sg13g2_FILL8
XSTDFILL15_2080 VDD VSS sg13g2_FILL8
XSTDFILL15_2088 VDD VSS sg13g2_FILL8
XSTDFILL15_2096 VDD VSS sg13g2_FILL8
XSTDFILL15_2104 VDD VSS sg13g2_FILL8
XSTDFILL15_2112 VDD VSS sg13g2_FILL8
XSTDFILL15_2120 VDD VSS sg13g2_FILL8
XSTDFILL15_2128 VDD VSS sg13g2_FILL8
XSTDFILL15_2136 VDD VSS sg13g2_FILL8
XSTDFILL15_2144 VDD VSS sg13g2_FILL8
XSTDFILL15_2152 VDD VSS sg13g2_FILL8
XSTDFILL15_2160 VDD VSS sg13g2_FILL8
XSTDFILL15_2168 VDD VSS sg13g2_FILL4
XSTDFILL16_0 VDD VSS sg13g2_FILL8
XSTDFILL16_8 VDD VSS sg13g2_FILL8
XSTDFILL16_16 VDD VSS sg13g2_FILL8
XSTDFILL16_24 VDD VSS sg13g2_FILL8
XSTDFILL16_32 VDD VSS sg13g2_FILL8
XSTDFILL16_40 VDD VSS sg13g2_FILL8
XSTDFILL16_48 VDD VSS sg13g2_FILL8
XSTDFILL16_56 VDD VSS sg13g2_FILL8
XSTDFILL16_64 VDD VSS sg13g2_FILL8
XSTDFILL16_72 VDD VSS sg13g2_FILL8
XSTDFILL16_80 VDD VSS sg13g2_FILL8
XSTDFILL16_88 VDD VSS sg13g2_FILL8
XSTDFILL16_96 VDD VSS sg13g2_FILL8
XSTDFILL16_104 VDD VSS sg13g2_FILL1
XSTDFILL16_1880 VDD VSS sg13g2_FILL8
XSTDFILL16_1888 VDD VSS sg13g2_FILL8
XSTDFILL16_1896 VDD VSS sg13g2_FILL8
XSTDFILL16_1904 VDD VSS sg13g2_FILL8
XSTDFILL16_1912 VDD VSS sg13g2_FILL8
XSTDFILL16_1920 VDD VSS sg13g2_FILL8
XSTDFILL16_1928 VDD VSS sg13g2_FILL8
XSTDFILL16_1936 VDD VSS sg13g2_FILL8
XSTDFILL16_1944 VDD VSS sg13g2_FILL8
XSTDFILL16_1952 VDD VSS sg13g2_FILL8
XSTDFILL16_1960 VDD VSS sg13g2_FILL8
XSTDFILL16_1968 VDD VSS sg13g2_FILL8
XSTDFILL16_1976 VDD VSS sg13g2_FILL8
XSTDFILL16_1984 VDD VSS sg13g2_FILL8
XSTDFILL16_1992 VDD VSS sg13g2_FILL8
XSTDFILL16_2000 VDD VSS sg13g2_FILL8
XSTDFILL16_2008 VDD VSS sg13g2_FILL8
XSTDFILL16_2016 VDD VSS sg13g2_FILL8
XSTDFILL16_2024 VDD VSS sg13g2_FILL8
XSTDFILL16_2032 VDD VSS sg13g2_FILL8
XSTDFILL16_2040 VDD VSS sg13g2_FILL8
XSTDFILL16_2048 VDD VSS sg13g2_FILL8
XSTDFILL16_2056 VDD VSS sg13g2_FILL8
XSTDFILL16_2064 VDD VSS sg13g2_FILL8
XSTDFILL16_2072 VDD VSS sg13g2_FILL8
XSTDFILL16_2080 VDD VSS sg13g2_FILL8
XSTDFILL16_2088 VDD VSS sg13g2_FILL8
XSTDFILL16_2096 VDD VSS sg13g2_FILL8
XSTDFILL16_2104 VDD VSS sg13g2_FILL8
XSTDFILL16_2112 VDD VSS sg13g2_FILL8
XSTDFILL16_2120 VDD VSS sg13g2_FILL8
XSTDFILL16_2128 VDD VSS sg13g2_FILL8
XSTDFILL16_2136 VDD VSS sg13g2_FILL8
XSTDFILL16_2144 VDD VSS sg13g2_FILL8
XSTDFILL16_2152 VDD VSS sg13g2_FILL8
XSTDFILL16_2160 VDD VSS sg13g2_FILL8
XSTDFILL16_2168 VDD VSS sg13g2_FILL4
XSTDFILL17_0 VDD VSS sg13g2_FILL8
XSTDFILL17_8 VDD VSS sg13g2_FILL8
XSTDFILL17_16 VDD VSS sg13g2_FILL8
XSTDFILL17_24 VDD VSS sg13g2_FILL8
XSTDFILL17_32 VDD VSS sg13g2_FILL8
XSTDFILL17_40 VDD VSS sg13g2_FILL8
XSTDFILL17_48 VDD VSS sg13g2_FILL8
XSTDFILL17_56 VDD VSS sg13g2_FILL8
XSTDFILL17_64 VDD VSS sg13g2_FILL8
XSTDFILL17_72 VDD VSS sg13g2_FILL8
XSTDFILL17_80 VDD VSS sg13g2_FILL8
XSTDFILL17_88 VDD VSS sg13g2_FILL8
XSTDFILL17_96 VDD VSS sg13g2_FILL8
XSTDFILL17_104 VDD VSS sg13g2_FILL1
XSTDFILL17_1880 VDD VSS sg13g2_FILL8
XSTDFILL17_1888 VDD VSS sg13g2_FILL8
XSTDFILL17_1896 VDD VSS sg13g2_FILL8
XSTDFILL17_1904 VDD VSS sg13g2_FILL8
XSTDFILL17_1912 VDD VSS sg13g2_FILL8
XSTDFILL17_1920 VDD VSS sg13g2_FILL8
XSTDFILL17_1928 VDD VSS sg13g2_FILL8
XSTDFILL17_1936 VDD VSS sg13g2_FILL8
XSTDFILL17_1944 VDD VSS sg13g2_FILL8
XSTDFILL17_1952 VDD VSS sg13g2_FILL8
XSTDFILL17_1960 VDD VSS sg13g2_FILL8
XSTDFILL17_1968 VDD VSS sg13g2_FILL8
XSTDFILL17_1976 VDD VSS sg13g2_FILL8
XSTDFILL17_1984 VDD VSS sg13g2_FILL8
XSTDFILL17_1992 VDD VSS sg13g2_FILL8
XSTDFILL17_2000 VDD VSS sg13g2_FILL8
XSTDFILL17_2008 VDD VSS sg13g2_FILL8
XSTDFILL17_2016 VDD VSS sg13g2_FILL8
XSTDFILL17_2024 VDD VSS sg13g2_FILL8
XSTDFILL17_2032 VDD VSS sg13g2_FILL8
XSTDFILL17_2040 VDD VSS sg13g2_FILL8
XSTDFILL17_2048 VDD VSS sg13g2_FILL8
XSTDFILL17_2056 VDD VSS sg13g2_FILL8
XSTDFILL17_2064 VDD VSS sg13g2_FILL8
XSTDFILL17_2072 VDD VSS sg13g2_FILL8
XSTDFILL17_2080 VDD VSS sg13g2_FILL8
XSTDFILL17_2088 VDD VSS sg13g2_FILL8
XSTDFILL17_2096 VDD VSS sg13g2_FILL8
XSTDFILL17_2104 VDD VSS sg13g2_FILL8
XSTDFILL17_2112 VDD VSS sg13g2_FILL8
XSTDFILL17_2120 VDD VSS sg13g2_FILL8
XSTDFILL17_2128 VDD VSS sg13g2_FILL8
XSTDFILL17_2136 VDD VSS sg13g2_FILL8
XSTDFILL17_2144 VDD VSS sg13g2_FILL8
XSTDFILL17_2152 VDD VSS sg13g2_FILL8
XSTDFILL17_2160 VDD VSS sg13g2_FILL8
XSTDFILL17_2168 VDD VSS sg13g2_FILL4
XSTDFILL18_0 VDD VSS sg13g2_FILL8
XSTDFILL18_8 VDD VSS sg13g2_FILL8
XSTDFILL18_16 VDD VSS sg13g2_FILL8
XSTDFILL18_24 VDD VSS sg13g2_FILL8
XSTDFILL18_32 VDD VSS sg13g2_FILL8
XSTDFILL18_40 VDD VSS sg13g2_FILL8
XSTDFILL18_48 VDD VSS sg13g2_FILL8
XSTDFILL18_56 VDD VSS sg13g2_FILL8
XSTDFILL18_64 VDD VSS sg13g2_FILL8
XSTDFILL18_72 VDD VSS sg13g2_FILL8
XSTDFILL18_80 VDD VSS sg13g2_FILL8
XSTDFILL18_88 VDD VSS sg13g2_FILL8
XSTDFILL18_96 VDD VSS sg13g2_FILL8
XSTDFILL18_104 VDD VSS sg13g2_FILL1
XSTDFILL18_1880 VDD VSS sg13g2_FILL8
XSTDFILL18_1888 VDD VSS sg13g2_FILL8
XSTDFILL18_1896 VDD VSS sg13g2_FILL8
XSTDFILL18_1904 VDD VSS sg13g2_FILL8
XSTDFILL18_1912 VDD VSS sg13g2_FILL8
XSTDFILL18_1920 VDD VSS sg13g2_FILL8
XSTDFILL18_1928 VDD VSS sg13g2_FILL8
XSTDFILL18_1936 VDD VSS sg13g2_FILL8
XSTDFILL18_1944 VDD VSS sg13g2_FILL8
XSTDFILL18_1952 VDD VSS sg13g2_FILL8
XSTDFILL18_1960 VDD VSS sg13g2_FILL8
XSTDFILL18_1968 VDD VSS sg13g2_FILL8
XSTDFILL18_1976 VDD VSS sg13g2_FILL8
XSTDFILL18_1984 VDD VSS sg13g2_FILL8
XSTDFILL18_1992 VDD VSS sg13g2_FILL8
XSTDFILL18_2000 VDD VSS sg13g2_FILL8
XSTDFILL18_2008 VDD VSS sg13g2_FILL8
XSTDFILL18_2016 VDD VSS sg13g2_FILL8
XSTDFILL18_2024 VDD VSS sg13g2_FILL8
XSTDFILL18_2032 VDD VSS sg13g2_FILL8
XSTDFILL18_2040 VDD VSS sg13g2_FILL8
XSTDFILL18_2048 VDD VSS sg13g2_FILL8
XSTDFILL18_2056 VDD VSS sg13g2_FILL8
XSTDFILL18_2064 VDD VSS sg13g2_FILL8
XSTDFILL18_2072 VDD VSS sg13g2_FILL8
XSTDFILL18_2080 VDD VSS sg13g2_FILL8
XSTDFILL18_2088 VDD VSS sg13g2_FILL8
XSTDFILL18_2096 VDD VSS sg13g2_FILL8
XSTDFILL18_2104 VDD VSS sg13g2_FILL8
XSTDFILL18_2112 VDD VSS sg13g2_FILL8
XSTDFILL18_2120 VDD VSS sg13g2_FILL8
XSTDFILL18_2128 VDD VSS sg13g2_FILL8
XSTDFILL18_2136 VDD VSS sg13g2_FILL8
XSTDFILL18_2144 VDD VSS sg13g2_FILL8
XSTDFILL18_2152 VDD VSS sg13g2_FILL8
XSTDFILL18_2160 VDD VSS sg13g2_FILL8
XSTDFILL18_2168 VDD VSS sg13g2_FILL4
XSTDFILL19_0 VDD VSS sg13g2_FILL8
XSTDFILL19_8 VDD VSS sg13g2_FILL8
XSTDFILL19_16 VDD VSS sg13g2_FILL8
XSTDFILL19_24 VDD VSS sg13g2_FILL8
XSTDFILL19_32 VDD VSS sg13g2_FILL8
XSTDFILL19_40 VDD VSS sg13g2_FILL8
XSTDFILL19_48 VDD VSS sg13g2_FILL8
XSTDFILL19_56 VDD VSS sg13g2_FILL8
XSTDFILL19_64 VDD VSS sg13g2_FILL8
XSTDFILL19_72 VDD VSS sg13g2_FILL8
XSTDFILL19_80 VDD VSS sg13g2_FILL8
XSTDFILL19_88 VDD VSS sg13g2_FILL8
XSTDFILL19_96 VDD VSS sg13g2_FILL8
XSTDFILL19_104 VDD VSS sg13g2_FILL1
XSTDFILL19_1880 VDD VSS sg13g2_FILL8
XSTDFILL19_1888 VDD VSS sg13g2_FILL8
XSTDFILL19_1896 VDD VSS sg13g2_FILL8
XSTDFILL19_1904 VDD VSS sg13g2_FILL8
XSTDFILL19_1912 VDD VSS sg13g2_FILL8
XSTDFILL19_1920 VDD VSS sg13g2_FILL8
XSTDFILL19_1928 VDD VSS sg13g2_FILL8
XSTDFILL19_1936 VDD VSS sg13g2_FILL8
XSTDFILL19_1944 VDD VSS sg13g2_FILL8
XSTDFILL19_1952 VDD VSS sg13g2_FILL8
XSTDFILL19_1960 VDD VSS sg13g2_FILL8
XSTDFILL19_1968 VDD VSS sg13g2_FILL8
XSTDFILL19_1976 VDD VSS sg13g2_FILL8
XSTDFILL19_1984 VDD VSS sg13g2_FILL8
XSTDFILL19_1992 VDD VSS sg13g2_FILL8
XSTDFILL19_2000 VDD VSS sg13g2_FILL8
XSTDFILL19_2008 VDD VSS sg13g2_FILL8
XSTDFILL19_2016 VDD VSS sg13g2_FILL8
XSTDFILL19_2024 VDD VSS sg13g2_FILL8
XSTDFILL19_2032 VDD VSS sg13g2_FILL8
XSTDFILL19_2040 VDD VSS sg13g2_FILL8
XSTDFILL19_2048 VDD VSS sg13g2_FILL8
XSTDFILL19_2056 VDD VSS sg13g2_FILL8
XSTDFILL19_2064 VDD VSS sg13g2_FILL8
XSTDFILL19_2072 VDD VSS sg13g2_FILL8
XSTDFILL19_2080 VDD VSS sg13g2_FILL8
XSTDFILL19_2088 VDD VSS sg13g2_FILL8
XSTDFILL19_2096 VDD VSS sg13g2_FILL8
XSTDFILL19_2104 VDD VSS sg13g2_FILL8
XSTDFILL19_2112 VDD VSS sg13g2_FILL8
XSTDFILL19_2120 VDD VSS sg13g2_FILL8
XSTDFILL19_2128 VDD VSS sg13g2_FILL8
XSTDFILL19_2136 VDD VSS sg13g2_FILL8
XSTDFILL19_2144 VDD VSS sg13g2_FILL8
XSTDFILL19_2152 VDD VSS sg13g2_FILL8
XSTDFILL19_2160 VDD VSS sg13g2_FILL8
XSTDFILL19_2168 VDD VSS sg13g2_FILL4
XSTDFILL20_0 VDD VSS sg13g2_FILL8
XSTDFILL20_8 VDD VSS sg13g2_FILL8
XSTDFILL20_16 VDD VSS sg13g2_FILL8
XSTDFILL20_24 VDD VSS sg13g2_FILL8
XSTDFILL20_32 VDD VSS sg13g2_FILL8
XSTDFILL20_40 VDD VSS sg13g2_FILL8
XSTDFILL20_48 VDD VSS sg13g2_FILL8
XSTDFILL20_56 VDD VSS sg13g2_FILL8
XSTDFILL20_64 VDD VSS sg13g2_FILL8
XSTDFILL20_72 VDD VSS sg13g2_FILL8
XSTDFILL20_80 VDD VSS sg13g2_FILL8
XSTDFILL20_88 VDD VSS sg13g2_FILL8
XSTDFILL20_96 VDD VSS sg13g2_FILL8
XSTDFILL20_104 VDD VSS sg13g2_FILL1
XSTDFILL20_1880 VDD VSS sg13g2_FILL8
XSTDFILL20_1888 VDD VSS sg13g2_FILL8
XSTDFILL20_1896 VDD VSS sg13g2_FILL8
XSTDFILL20_1904 VDD VSS sg13g2_FILL8
XSTDFILL20_1912 VDD VSS sg13g2_FILL8
XSTDFILL20_1920 VDD VSS sg13g2_FILL8
XSTDFILL20_1928 VDD VSS sg13g2_FILL8
XSTDFILL20_1936 VDD VSS sg13g2_FILL8
XSTDFILL20_1944 VDD VSS sg13g2_FILL8
XSTDFILL20_1952 VDD VSS sg13g2_FILL8
XSTDFILL20_1960 VDD VSS sg13g2_FILL8
XSTDFILL20_1968 VDD VSS sg13g2_FILL8
XSTDFILL20_1976 VDD VSS sg13g2_FILL8
XSTDFILL20_1984 VDD VSS sg13g2_FILL8
XSTDFILL20_1992 VDD VSS sg13g2_FILL8
XSTDFILL20_2000 VDD VSS sg13g2_FILL8
XSTDFILL20_2008 VDD VSS sg13g2_FILL8
XSTDFILL20_2016 VDD VSS sg13g2_FILL8
XSTDFILL20_2024 VDD VSS sg13g2_FILL8
XSTDFILL20_2032 VDD VSS sg13g2_FILL8
XSTDFILL20_2040 VDD VSS sg13g2_FILL8
XSTDFILL20_2048 VDD VSS sg13g2_FILL8
XSTDFILL20_2056 VDD VSS sg13g2_FILL8
XSTDFILL20_2064 VDD VSS sg13g2_FILL8
XSTDFILL20_2072 VDD VSS sg13g2_FILL8
XSTDFILL20_2080 VDD VSS sg13g2_FILL8
XSTDFILL20_2088 VDD VSS sg13g2_FILL8
XSTDFILL20_2096 VDD VSS sg13g2_FILL8
XSTDFILL20_2104 VDD VSS sg13g2_FILL8
XSTDFILL20_2112 VDD VSS sg13g2_FILL8
XSTDFILL20_2120 VDD VSS sg13g2_FILL8
XSTDFILL20_2128 VDD VSS sg13g2_FILL8
XSTDFILL20_2136 VDD VSS sg13g2_FILL8
XSTDFILL20_2144 VDD VSS sg13g2_FILL8
XSTDFILL20_2152 VDD VSS sg13g2_FILL8
XSTDFILL20_2160 VDD VSS sg13g2_FILL8
XSTDFILL20_2168 VDD VSS sg13g2_FILL4
XSTDFILL21_0 VDD VSS sg13g2_FILL8
XSTDFILL21_8 VDD VSS sg13g2_FILL8
XSTDFILL21_16 VDD VSS sg13g2_FILL8
XSTDFILL21_24 VDD VSS sg13g2_FILL8
XSTDFILL21_32 VDD VSS sg13g2_FILL8
XSTDFILL21_40 VDD VSS sg13g2_FILL8
XSTDFILL21_48 VDD VSS sg13g2_FILL8
XSTDFILL21_56 VDD VSS sg13g2_FILL8
XSTDFILL21_64 VDD VSS sg13g2_FILL8
XSTDFILL21_72 VDD VSS sg13g2_FILL8
XSTDFILL21_80 VDD VSS sg13g2_FILL8
XSTDFILL21_88 VDD VSS sg13g2_FILL8
XSTDFILL21_96 VDD VSS sg13g2_FILL8
XSTDFILL21_104 VDD VSS sg13g2_FILL1
XSTDFILL21_1880 VDD VSS sg13g2_FILL8
XSTDFILL21_1888 VDD VSS sg13g2_FILL8
XSTDFILL21_1896 VDD VSS sg13g2_FILL8
XSTDFILL21_1904 VDD VSS sg13g2_FILL8
XSTDFILL21_1912 VDD VSS sg13g2_FILL8
XSTDFILL21_1920 VDD VSS sg13g2_FILL8
XSTDFILL21_1928 VDD VSS sg13g2_FILL8
XSTDFILL21_1936 VDD VSS sg13g2_FILL8
XSTDFILL21_1944 VDD VSS sg13g2_FILL8
XSTDFILL21_1952 VDD VSS sg13g2_FILL8
XSTDFILL21_1960 VDD VSS sg13g2_FILL8
XSTDFILL21_1968 VDD VSS sg13g2_FILL8
XSTDFILL21_1976 VDD VSS sg13g2_FILL8
XSTDFILL21_1984 VDD VSS sg13g2_FILL8
XSTDFILL21_1992 VDD VSS sg13g2_FILL8
XSTDFILL21_2000 VDD VSS sg13g2_FILL8
XSTDFILL21_2008 VDD VSS sg13g2_FILL8
XSTDFILL21_2016 VDD VSS sg13g2_FILL8
XSTDFILL21_2024 VDD VSS sg13g2_FILL8
XSTDFILL21_2032 VDD VSS sg13g2_FILL8
XSTDFILL21_2040 VDD VSS sg13g2_FILL8
XSTDFILL21_2048 VDD VSS sg13g2_FILL8
XSTDFILL21_2056 VDD VSS sg13g2_FILL8
XSTDFILL21_2064 VDD VSS sg13g2_FILL8
XSTDFILL21_2072 VDD VSS sg13g2_FILL8
XSTDFILL21_2080 VDD VSS sg13g2_FILL8
XSTDFILL21_2088 VDD VSS sg13g2_FILL8
XSTDFILL21_2096 VDD VSS sg13g2_FILL8
XSTDFILL21_2104 VDD VSS sg13g2_FILL8
XSTDFILL21_2112 VDD VSS sg13g2_FILL8
XSTDFILL21_2120 VDD VSS sg13g2_FILL8
XSTDFILL21_2128 VDD VSS sg13g2_FILL8
XSTDFILL21_2136 VDD VSS sg13g2_FILL8
XSTDFILL21_2144 VDD VSS sg13g2_FILL8
XSTDFILL21_2152 VDD VSS sg13g2_FILL8
XSTDFILL21_2160 VDD VSS sg13g2_FILL8
XSTDFILL21_2168 VDD VSS sg13g2_FILL4
XSTDFILL22_0 VDD VSS sg13g2_FILL8
XSTDFILL22_8 VDD VSS sg13g2_FILL8
XSTDFILL22_16 VDD VSS sg13g2_FILL8
XSTDFILL22_24 VDD VSS sg13g2_FILL8
XSTDFILL22_32 VDD VSS sg13g2_FILL8
XSTDFILL22_40 VDD VSS sg13g2_FILL8
XSTDFILL22_48 VDD VSS sg13g2_FILL8
XSTDFILL22_56 VDD VSS sg13g2_FILL8
XSTDFILL22_64 VDD VSS sg13g2_FILL8
XSTDFILL22_72 VDD VSS sg13g2_FILL8
XSTDFILL22_80 VDD VSS sg13g2_FILL8
XSTDFILL22_88 VDD VSS sg13g2_FILL8
XSTDFILL22_96 VDD VSS sg13g2_FILL8
XSTDFILL22_104 VDD VSS sg13g2_FILL1
XSTDFILL22_1880 VDD VSS sg13g2_FILL8
XSTDFILL22_1888 VDD VSS sg13g2_FILL8
XSTDFILL22_1896 VDD VSS sg13g2_FILL8
XSTDFILL22_1904 VDD VSS sg13g2_FILL8
XSTDFILL22_1912 VDD VSS sg13g2_FILL8
XSTDFILL22_1920 VDD VSS sg13g2_FILL8
XSTDFILL22_1928 VDD VSS sg13g2_FILL8
XSTDFILL22_1936 VDD VSS sg13g2_FILL8
XSTDFILL22_1944 VDD VSS sg13g2_FILL8
XSTDFILL22_1952 VDD VSS sg13g2_FILL8
XSTDFILL22_1960 VDD VSS sg13g2_FILL8
XSTDFILL22_1968 VDD VSS sg13g2_FILL8
XSTDFILL22_1976 VDD VSS sg13g2_FILL8
XSTDFILL22_1984 VDD VSS sg13g2_FILL8
XSTDFILL22_1992 VDD VSS sg13g2_FILL8
XSTDFILL22_2000 VDD VSS sg13g2_FILL8
XSTDFILL22_2008 VDD VSS sg13g2_FILL8
XSTDFILL22_2016 VDD VSS sg13g2_FILL8
XSTDFILL22_2024 VDD VSS sg13g2_FILL8
XSTDFILL22_2032 VDD VSS sg13g2_FILL8
XSTDFILL22_2040 VDD VSS sg13g2_FILL8
XSTDFILL22_2048 VDD VSS sg13g2_FILL8
XSTDFILL22_2056 VDD VSS sg13g2_FILL8
XSTDFILL22_2064 VDD VSS sg13g2_FILL8
XSTDFILL22_2072 VDD VSS sg13g2_FILL8
XSTDFILL22_2080 VDD VSS sg13g2_FILL8
XSTDFILL22_2088 VDD VSS sg13g2_FILL8
XSTDFILL22_2096 VDD VSS sg13g2_FILL8
XSTDFILL22_2104 VDD VSS sg13g2_FILL8
XSTDFILL22_2112 VDD VSS sg13g2_FILL8
XSTDFILL22_2120 VDD VSS sg13g2_FILL8
XSTDFILL22_2128 VDD VSS sg13g2_FILL8
XSTDFILL22_2136 VDD VSS sg13g2_FILL8
XSTDFILL22_2144 VDD VSS sg13g2_FILL8
XSTDFILL22_2152 VDD VSS sg13g2_FILL8
XSTDFILL22_2160 VDD VSS sg13g2_FILL8
XSTDFILL22_2168 VDD VSS sg13g2_FILL4
XSTDFILL23_0 VDD VSS sg13g2_FILL8
XSTDFILL23_8 VDD VSS sg13g2_FILL8
XSTDFILL23_16 VDD VSS sg13g2_FILL8
XSTDFILL23_24 VDD VSS sg13g2_FILL8
XSTDFILL23_32 VDD VSS sg13g2_FILL8
XSTDFILL23_40 VDD VSS sg13g2_FILL8
XSTDFILL23_48 VDD VSS sg13g2_FILL8
XSTDFILL23_56 VDD VSS sg13g2_FILL8
XSTDFILL23_64 VDD VSS sg13g2_FILL8
XSTDFILL23_72 VDD VSS sg13g2_FILL8
XSTDFILL23_80 VDD VSS sg13g2_FILL8
XSTDFILL23_88 VDD VSS sg13g2_FILL8
XSTDFILL23_96 VDD VSS sg13g2_FILL8
XSTDFILL23_104 VDD VSS sg13g2_FILL1
XSTDFILL23_1880 VDD VSS sg13g2_FILL8
XSTDFILL23_1888 VDD VSS sg13g2_FILL8
XSTDFILL23_1896 VDD VSS sg13g2_FILL8
XSTDFILL23_1904 VDD VSS sg13g2_FILL8
XSTDFILL23_1912 VDD VSS sg13g2_FILL8
XSTDFILL23_1920 VDD VSS sg13g2_FILL8
XSTDFILL23_1928 VDD VSS sg13g2_FILL8
XSTDFILL23_1936 VDD VSS sg13g2_FILL8
XSTDFILL23_1944 VDD VSS sg13g2_FILL8
XSTDFILL23_1952 VDD VSS sg13g2_FILL8
XSTDFILL23_1960 VDD VSS sg13g2_FILL8
XSTDFILL23_1968 VDD VSS sg13g2_FILL8
XSTDFILL23_1976 VDD VSS sg13g2_FILL8
XSTDFILL23_1984 VDD VSS sg13g2_FILL8
XSTDFILL23_1992 VDD VSS sg13g2_FILL8
XSTDFILL23_2000 VDD VSS sg13g2_FILL8
XSTDFILL23_2008 VDD VSS sg13g2_FILL8
XSTDFILL23_2016 VDD VSS sg13g2_FILL8
XSTDFILL23_2024 VDD VSS sg13g2_FILL8
XSTDFILL23_2032 VDD VSS sg13g2_FILL8
XSTDFILL23_2040 VDD VSS sg13g2_FILL8
XSTDFILL23_2048 VDD VSS sg13g2_FILL8
XSTDFILL23_2056 VDD VSS sg13g2_FILL8
XSTDFILL23_2064 VDD VSS sg13g2_FILL8
XSTDFILL23_2072 VDD VSS sg13g2_FILL8
XSTDFILL23_2080 VDD VSS sg13g2_FILL8
XSTDFILL23_2088 VDD VSS sg13g2_FILL8
XSTDFILL23_2096 VDD VSS sg13g2_FILL8
XSTDFILL23_2104 VDD VSS sg13g2_FILL8
XSTDFILL23_2112 VDD VSS sg13g2_FILL8
XSTDFILL23_2120 VDD VSS sg13g2_FILL8
XSTDFILL23_2128 VDD VSS sg13g2_FILL8
XSTDFILL23_2136 VDD VSS sg13g2_FILL8
XSTDFILL23_2144 VDD VSS sg13g2_FILL8
XSTDFILL23_2152 VDD VSS sg13g2_FILL8
XSTDFILL23_2160 VDD VSS sg13g2_FILL8
XSTDFILL23_2168 VDD VSS sg13g2_FILL4
XSTDFILL24_0 VDD VSS sg13g2_FILL8
XSTDFILL24_8 VDD VSS sg13g2_FILL8
XSTDFILL24_16 VDD VSS sg13g2_FILL8
XSTDFILL24_24 VDD VSS sg13g2_FILL8
XSTDFILL24_32 VDD VSS sg13g2_FILL8
XSTDFILL24_40 VDD VSS sg13g2_FILL8
XSTDFILL24_48 VDD VSS sg13g2_FILL8
XSTDFILL24_56 VDD VSS sg13g2_FILL8
XSTDFILL24_64 VDD VSS sg13g2_FILL8
XSTDFILL24_72 VDD VSS sg13g2_FILL8
XSTDFILL24_80 VDD VSS sg13g2_FILL8
XSTDFILL24_88 VDD VSS sg13g2_FILL8
XSTDFILL24_96 VDD VSS sg13g2_FILL8
XSTDFILL24_104 VDD VSS sg13g2_FILL1
XSTDFILL24_1880 VDD VSS sg13g2_FILL8
XSTDFILL24_1888 VDD VSS sg13g2_FILL8
XSTDFILL24_1896 VDD VSS sg13g2_FILL8
XSTDFILL24_1904 VDD VSS sg13g2_FILL8
XSTDFILL24_1912 VDD VSS sg13g2_FILL8
XSTDFILL24_1920 VDD VSS sg13g2_FILL8
XSTDFILL24_1928 VDD VSS sg13g2_FILL8
XSTDFILL24_1936 VDD VSS sg13g2_FILL8
XSTDFILL24_1944 VDD VSS sg13g2_FILL8
XSTDFILL24_1952 VDD VSS sg13g2_FILL8
XSTDFILL24_1960 VDD VSS sg13g2_FILL8
XSTDFILL24_1968 VDD VSS sg13g2_FILL8
XSTDFILL24_1976 VDD VSS sg13g2_FILL8
XSTDFILL24_1984 VDD VSS sg13g2_FILL8
XSTDFILL24_1992 VDD VSS sg13g2_FILL8
XSTDFILL24_2000 VDD VSS sg13g2_FILL8
XSTDFILL24_2008 VDD VSS sg13g2_FILL8
XSTDFILL24_2016 VDD VSS sg13g2_FILL8
XSTDFILL24_2024 VDD VSS sg13g2_FILL8
XSTDFILL24_2032 VDD VSS sg13g2_FILL8
XSTDFILL24_2040 VDD VSS sg13g2_FILL8
XSTDFILL24_2048 VDD VSS sg13g2_FILL8
XSTDFILL24_2056 VDD VSS sg13g2_FILL8
XSTDFILL24_2064 VDD VSS sg13g2_FILL8
XSTDFILL24_2072 VDD VSS sg13g2_FILL8
XSTDFILL24_2080 VDD VSS sg13g2_FILL8
XSTDFILL24_2088 VDD VSS sg13g2_FILL8
XSTDFILL24_2096 VDD VSS sg13g2_FILL8
XSTDFILL24_2104 VDD VSS sg13g2_FILL8
XSTDFILL24_2112 VDD VSS sg13g2_FILL8
XSTDFILL24_2120 VDD VSS sg13g2_FILL8
XSTDFILL24_2128 VDD VSS sg13g2_FILL8
XSTDFILL24_2136 VDD VSS sg13g2_FILL8
XSTDFILL24_2144 VDD VSS sg13g2_FILL8
XSTDFILL24_2152 VDD VSS sg13g2_FILL8
XSTDFILL24_2160 VDD VSS sg13g2_FILL8
XSTDFILL24_2168 VDD VSS sg13g2_FILL4
XSTDFILL25_0 VDD VSS sg13g2_FILL8
XSTDFILL25_8 VDD VSS sg13g2_FILL8
XSTDFILL25_16 VDD VSS sg13g2_FILL8
XSTDFILL25_24 VDD VSS sg13g2_FILL8
XSTDFILL25_32 VDD VSS sg13g2_FILL8
XSTDFILL25_40 VDD VSS sg13g2_FILL8
XSTDFILL25_48 VDD VSS sg13g2_FILL8
XSTDFILL25_56 VDD VSS sg13g2_FILL8
XSTDFILL25_64 VDD VSS sg13g2_FILL8
XSTDFILL25_72 VDD VSS sg13g2_FILL8
XSTDFILL25_80 VDD VSS sg13g2_FILL8
XSTDFILL25_88 VDD VSS sg13g2_FILL8
XSTDFILL25_96 VDD VSS sg13g2_FILL8
XSTDFILL25_104 VDD VSS sg13g2_FILL1
XSTDFILL25_1880 VDD VSS sg13g2_FILL8
XSTDFILL25_1888 VDD VSS sg13g2_FILL8
XSTDFILL25_1896 VDD VSS sg13g2_FILL8
XSTDFILL25_1904 VDD VSS sg13g2_FILL8
XSTDFILL25_1912 VDD VSS sg13g2_FILL8
XSTDFILL25_1920 VDD VSS sg13g2_FILL8
XSTDFILL25_1928 VDD VSS sg13g2_FILL8
XSTDFILL25_1936 VDD VSS sg13g2_FILL8
XSTDFILL25_1944 VDD VSS sg13g2_FILL8
XSTDFILL25_1952 VDD VSS sg13g2_FILL8
XSTDFILL25_1960 VDD VSS sg13g2_FILL8
XSTDFILL25_1968 VDD VSS sg13g2_FILL8
XSTDFILL25_1976 VDD VSS sg13g2_FILL8
XSTDFILL25_1984 VDD VSS sg13g2_FILL8
XSTDFILL25_1992 VDD VSS sg13g2_FILL8
XSTDFILL25_2000 VDD VSS sg13g2_FILL8
XSTDFILL25_2008 VDD VSS sg13g2_FILL8
XSTDFILL25_2016 VDD VSS sg13g2_FILL8
XSTDFILL25_2024 VDD VSS sg13g2_FILL8
XSTDFILL25_2032 VDD VSS sg13g2_FILL8
XSTDFILL25_2040 VDD VSS sg13g2_FILL8
XSTDFILL25_2048 VDD VSS sg13g2_FILL8
XSTDFILL25_2056 VDD VSS sg13g2_FILL8
XSTDFILL25_2064 VDD VSS sg13g2_FILL8
XSTDFILL25_2072 VDD VSS sg13g2_FILL8
XSTDFILL25_2080 VDD VSS sg13g2_FILL8
XSTDFILL25_2088 VDD VSS sg13g2_FILL8
XSTDFILL25_2096 VDD VSS sg13g2_FILL8
XSTDFILL25_2104 VDD VSS sg13g2_FILL8
XSTDFILL25_2112 VDD VSS sg13g2_FILL8
XSTDFILL25_2120 VDD VSS sg13g2_FILL8
XSTDFILL25_2128 VDD VSS sg13g2_FILL8
XSTDFILL25_2136 VDD VSS sg13g2_FILL8
XSTDFILL25_2144 VDD VSS sg13g2_FILL8
XSTDFILL25_2152 VDD VSS sg13g2_FILL8
XSTDFILL25_2160 VDD VSS sg13g2_FILL8
XSTDFILL25_2168 VDD VSS sg13g2_FILL4
XSTDFILL26_0 VDD VSS sg13g2_FILL8
XSTDFILL26_8 VDD VSS sg13g2_FILL8
XSTDFILL26_16 VDD VSS sg13g2_FILL8
XSTDFILL26_24 VDD VSS sg13g2_FILL8
XSTDFILL26_32 VDD VSS sg13g2_FILL8
XSTDFILL26_40 VDD VSS sg13g2_FILL8
XSTDFILL26_48 VDD VSS sg13g2_FILL8
XSTDFILL26_56 VDD VSS sg13g2_FILL8
XSTDFILL26_64 VDD VSS sg13g2_FILL8
XSTDFILL26_72 VDD VSS sg13g2_FILL8
XSTDFILL26_80 VDD VSS sg13g2_FILL8
XSTDFILL26_88 VDD VSS sg13g2_FILL8
XSTDFILL26_96 VDD VSS sg13g2_FILL8
XSTDFILL26_104 VDD VSS sg13g2_FILL1
XSTDFILL26_1880 VDD VSS sg13g2_FILL8
XSTDFILL26_1888 VDD VSS sg13g2_FILL8
XSTDFILL26_1896 VDD VSS sg13g2_FILL8
XSTDFILL26_1904 VDD VSS sg13g2_FILL8
XSTDFILL26_1912 VDD VSS sg13g2_FILL8
XSTDFILL26_1920 VDD VSS sg13g2_FILL8
XSTDFILL26_1928 VDD VSS sg13g2_FILL8
XSTDFILL26_1936 VDD VSS sg13g2_FILL8
XSTDFILL26_1944 VDD VSS sg13g2_FILL8
XSTDFILL26_1952 VDD VSS sg13g2_FILL8
XSTDFILL26_1960 VDD VSS sg13g2_FILL8
XSTDFILL26_1968 VDD VSS sg13g2_FILL8
XSTDFILL26_1976 VDD VSS sg13g2_FILL8
XSTDFILL26_1984 VDD VSS sg13g2_FILL8
XSTDFILL26_1992 VDD VSS sg13g2_FILL8
XSTDFILL26_2000 VDD VSS sg13g2_FILL8
XSTDFILL26_2008 VDD VSS sg13g2_FILL8
XSTDFILL26_2016 VDD VSS sg13g2_FILL8
XSTDFILL26_2024 VDD VSS sg13g2_FILL8
XSTDFILL26_2032 VDD VSS sg13g2_FILL8
XSTDFILL26_2040 VDD VSS sg13g2_FILL8
XSTDFILL26_2048 VDD VSS sg13g2_FILL8
XSTDFILL26_2056 VDD VSS sg13g2_FILL8
XSTDFILL26_2064 VDD VSS sg13g2_FILL8
XSTDFILL26_2072 VDD VSS sg13g2_FILL8
XSTDFILL26_2080 VDD VSS sg13g2_FILL8
XSTDFILL26_2088 VDD VSS sg13g2_FILL8
XSTDFILL26_2096 VDD VSS sg13g2_FILL8
XSTDFILL26_2104 VDD VSS sg13g2_FILL8
XSTDFILL26_2112 VDD VSS sg13g2_FILL8
XSTDFILL26_2120 VDD VSS sg13g2_FILL8
XSTDFILL26_2128 VDD VSS sg13g2_FILL8
XSTDFILL26_2136 VDD VSS sg13g2_FILL8
XSTDFILL26_2144 VDD VSS sg13g2_FILL8
XSTDFILL26_2152 VDD VSS sg13g2_FILL8
XSTDFILL26_2160 VDD VSS sg13g2_FILL8
XSTDFILL26_2168 VDD VSS sg13g2_FILL4
XSTDFILL27_0 VDD VSS sg13g2_FILL8
XSTDFILL27_8 VDD VSS sg13g2_FILL8
XSTDFILL27_16 VDD VSS sg13g2_FILL8
XSTDFILL27_24 VDD VSS sg13g2_FILL8
XSTDFILL27_32 VDD VSS sg13g2_FILL8
XSTDFILL27_40 VDD VSS sg13g2_FILL8
XSTDFILL27_48 VDD VSS sg13g2_FILL8
XSTDFILL27_56 VDD VSS sg13g2_FILL8
XSTDFILL27_64 VDD VSS sg13g2_FILL8
XSTDFILL27_72 VDD VSS sg13g2_FILL8
XSTDFILL27_80 VDD VSS sg13g2_FILL8
XSTDFILL27_88 VDD VSS sg13g2_FILL8
XSTDFILL27_96 VDD VSS sg13g2_FILL8
XSTDFILL27_104 VDD VSS sg13g2_FILL1
XSTDFILL27_1880 VDD VSS sg13g2_FILL8
XSTDFILL27_1888 VDD VSS sg13g2_FILL8
XSTDFILL27_1896 VDD VSS sg13g2_FILL8
XSTDFILL27_1904 VDD VSS sg13g2_FILL8
XSTDFILL27_1912 VDD VSS sg13g2_FILL8
XSTDFILL27_1920 VDD VSS sg13g2_FILL8
XSTDFILL27_1928 VDD VSS sg13g2_FILL8
XSTDFILL27_1936 VDD VSS sg13g2_FILL8
XSTDFILL27_1944 VDD VSS sg13g2_FILL8
XSTDFILL27_1952 VDD VSS sg13g2_FILL8
XSTDFILL27_1960 VDD VSS sg13g2_FILL8
XSTDFILL27_1968 VDD VSS sg13g2_FILL8
XSTDFILL27_1976 VDD VSS sg13g2_FILL8
XSTDFILL27_1984 VDD VSS sg13g2_FILL8
XSTDFILL27_1992 VDD VSS sg13g2_FILL8
XSTDFILL27_2000 VDD VSS sg13g2_FILL8
XSTDFILL27_2008 VDD VSS sg13g2_FILL8
XSTDFILL27_2016 VDD VSS sg13g2_FILL8
XSTDFILL27_2024 VDD VSS sg13g2_FILL8
XSTDFILL27_2032 VDD VSS sg13g2_FILL8
XSTDFILL27_2040 VDD VSS sg13g2_FILL8
XSTDFILL27_2048 VDD VSS sg13g2_FILL8
XSTDFILL27_2056 VDD VSS sg13g2_FILL8
XSTDFILL27_2064 VDD VSS sg13g2_FILL8
XSTDFILL27_2072 VDD VSS sg13g2_FILL8
XSTDFILL27_2080 VDD VSS sg13g2_FILL8
XSTDFILL27_2088 VDD VSS sg13g2_FILL8
XSTDFILL27_2096 VDD VSS sg13g2_FILL8
XSTDFILL27_2104 VDD VSS sg13g2_FILL8
XSTDFILL27_2112 VDD VSS sg13g2_FILL8
XSTDFILL27_2120 VDD VSS sg13g2_FILL8
XSTDFILL27_2128 VDD VSS sg13g2_FILL8
XSTDFILL27_2136 VDD VSS sg13g2_FILL8
XSTDFILL27_2144 VDD VSS sg13g2_FILL8
XSTDFILL27_2152 VDD VSS sg13g2_FILL8
XSTDFILL27_2160 VDD VSS sg13g2_FILL8
XSTDFILL27_2168 VDD VSS sg13g2_FILL4
XSTDFILL28_0 VDD VSS sg13g2_FILL8
XSTDFILL28_8 VDD VSS sg13g2_FILL8
XSTDFILL28_16 VDD VSS sg13g2_FILL8
XSTDFILL28_24 VDD VSS sg13g2_FILL8
XSTDFILL28_32 VDD VSS sg13g2_FILL8
XSTDFILL28_40 VDD VSS sg13g2_FILL8
XSTDFILL28_48 VDD VSS sg13g2_FILL8
XSTDFILL28_56 VDD VSS sg13g2_FILL8
XSTDFILL28_64 VDD VSS sg13g2_FILL8
XSTDFILL28_72 VDD VSS sg13g2_FILL8
XSTDFILL28_80 VDD VSS sg13g2_FILL8
XSTDFILL28_88 VDD VSS sg13g2_FILL8
XSTDFILL28_96 VDD VSS sg13g2_FILL8
XSTDFILL28_104 VDD VSS sg13g2_FILL1
XSTDFILL28_1880 VDD VSS sg13g2_FILL8
XSTDFILL28_1888 VDD VSS sg13g2_FILL8
XSTDFILL28_1896 VDD VSS sg13g2_FILL8
XSTDFILL28_1904 VDD VSS sg13g2_FILL8
XSTDFILL28_1912 VDD VSS sg13g2_FILL8
XSTDFILL28_1920 VDD VSS sg13g2_FILL8
XSTDFILL28_1928 VDD VSS sg13g2_FILL8
XSTDFILL28_1936 VDD VSS sg13g2_FILL8
XSTDFILL28_1944 VDD VSS sg13g2_FILL8
XSTDFILL28_1952 VDD VSS sg13g2_FILL8
XSTDFILL28_1960 VDD VSS sg13g2_FILL8
XSTDFILL28_1968 VDD VSS sg13g2_FILL8
XSTDFILL28_1976 VDD VSS sg13g2_FILL8
XSTDFILL28_1984 VDD VSS sg13g2_FILL8
XSTDFILL28_1992 VDD VSS sg13g2_FILL8
XSTDFILL28_2000 VDD VSS sg13g2_FILL8
XSTDFILL28_2008 VDD VSS sg13g2_FILL8
XSTDFILL28_2016 VDD VSS sg13g2_FILL8
XSTDFILL28_2024 VDD VSS sg13g2_FILL8
XSTDFILL28_2032 VDD VSS sg13g2_FILL8
XSTDFILL28_2040 VDD VSS sg13g2_FILL8
XSTDFILL28_2048 VDD VSS sg13g2_FILL8
XSTDFILL28_2056 VDD VSS sg13g2_FILL8
XSTDFILL28_2064 VDD VSS sg13g2_FILL8
XSTDFILL28_2072 VDD VSS sg13g2_FILL8
XSTDFILL28_2080 VDD VSS sg13g2_FILL8
XSTDFILL28_2088 VDD VSS sg13g2_FILL8
XSTDFILL28_2096 VDD VSS sg13g2_FILL8
XSTDFILL28_2104 VDD VSS sg13g2_FILL8
XSTDFILL28_2112 VDD VSS sg13g2_FILL8
XSTDFILL28_2120 VDD VSS sg13g2_FILL8
XSTDFILL28_2128 VDD VSS sg13g2_FILL8
XSTDFILL28_2136 VDD VSS sg13g2_FILL8
XSTDFILL28_2144 VDD VSS sg13g2_FILL8
XSTDFILL28_2152 VDD VSS sg13g2_FILL8
XSTDFILL28_2160 VDD VSS sg13g2_FILL8
XSTDFILL28_2168 VDD VSS sg13g2_FILL4
XSTDFILL29_0 VDD VSS sg13g2_FILL8
XSTDFILL29_8 VDD VSS sg13g2_FILL8
XSTDFILL29_16 VDD VSS sg13g2_FILL8
XSTDFILL29_24 VDD VSS sg13g2_FILL8
XSTDFILL29_32 VDD VSS sg13g2_FILL8
XSTDFILL29_40 VDD VSS sg13g2_FILL8
XSTDFILL29_48 VDD VSS sg13g2_FILL8
XSTDFILL29_56 VDD VSS sg13g2_FILL8
XSTDFILL29_64 VDD VSS sg13g2_FILL8
XSTDFILL29_72 VDD VSS sg13g2_FILL8
XSTDFILL29_80 VDD VSS sg13g2_FILL8
XSTDFILL29_88 VDD VSS sg13g2_FILL8
XSTDFILL29_96 VDD VSS sg13g2_FILL8
XSTDFILL29_104 VDD VSS sg13g2_FILL1
XSTDFILL29_1880 VDD VSS sg13g2_FILL8
XSTDFILL29_1888 VDD VSS sg13g2_FILL8
XSTDFILL29_1896 VDD VSS sg13g2_FILL8
XSTDFILL29_1904 VDD VSS sg13g2_FILL8
XSTDFILL29_1912 VDD VSS sg13g2_FILL8
XSTDFILL29_1920 VDD VSS sg13g2_FILL8
XSTDFILL29_1928 VDD VSS sg13g2_FILL8
XSTDFILL29_1936 VDD VSS sg13g2_FILL8
XSTDFILL29_1944 VDD VSS sg13g2_FILL8
XSTDFILL29_1952 VDD VSS sg13g2_FILL8
XSTDFILL29_1960 VDD VSS sg13g2_FILL8
XSTDFILL29_1968 VDD VSS sg13g2_FILL8
XSTDFILL29_1976 VDD VSS sg13g2_FILL8
XSTDFILL29_1984 VDD VSS sg13g2_FILL8
XSTDFILL29_1992 VDD VSS sg13g2_FILL8
XSTDFILL29_2000 VDD VSS sg13g2_FILL8
XSTDFILL29_2008 VDD VSS sg13g2_FILL8
XSTDFILL29_2016 VDD VSS sg13g2_FILL8
XSTDFILL29_2024 VDD VSS sg13g2_FILL8
XSTDFILL29_2032 VDD VSS sg13g2_FILL8
XSTDFILL29_2040 VDD VSS sg13g2_FILL8
XSTDFILL29_2048 VDD VSS sg13g2_FILL8
XSTDFILL29_2056 VDD VSS sg13g2_FILL8
XSTDFILL29_2064 VDD VSS sg13g2_FILL8
XSTDFILL29_2072 VDD VSS sg13g2_FILL8
XSTDFILL29_2080 VDD VSS sg13g2_FILL8
XSTDFILL29_2088 VDD VSS sg13g2_FILL8
XSTDFILL29_2096 VDD VSS sg13g2_FILL8
XSTDFILL29_2104 VDD VSS sg13g2_FILL8
XSTDFILL29_2112 VDD VSS sg13g2_FILL8
XSTDFILL29_2120 VDD VSS sg13g2_FILL8
XSTDFILL29_2128 VDD VSS sg13g2_FILL8
XSTDFILL29_2136 VDD VSS sg13g2_FILL8
XSTDFILL29_2144 VDD VSS sg13g2_FILL8
XSTDFILL29_2152 VDD VSS sg13g2_FILL8
XSTDFILL29_2160 VDD VSS sg13g2_FILL8
XSTDFILL29_2168 VDD VSS sg13g2_FILL4
XSTDFILL30_0 VDD VSS sg13g2_FILL8
XSTDFILL30_8 VDD VSS sg13g2_FILL8
XSTDFILL30_16 VDD VSS sg13g2_FILL8
XSTDFILL30_24 VDD VSS sg13g2_FILL8
XSTDFILL30_32 VDD VSS sg13g2_FILL8
XSTDFILL30_40 VDD VSS sg13g2_FILL8
XSTDFILL30_48 VDD VSS sg13g2_FILL8
XSTDFILL30_56 VDD VSS sg13g2_FILL8
XSTDFILL30_64 VDD VSS sg13g2_FILL8
XSTDFILL30_72 VDD VSS sg13g2_FILL8
XSTDFILL30_80 VDD VSS sg13g2_FILL8
XSTDFILL30_88 VDD VSS sg13g2_FILL8
XSTDFILL30_96 VDD VSS sg13g2_FILL8
XSTDFILL30_104 VDD VSS sg13g2_FILL1
XSTDFILL30_1880 VDD VSS sg13g2_FILL8
XSTDFILL30_1888 VDD VSS sg13g2_FILL8
XSTDFILL30_1896 VDD VSS sg13g2_FILL8
XSTDFILL30_1904 VDD VSS sg13g2_FILL8
XSTDFILL30_1912 VDD VSS sg13g2_FILL8
XSTDFILL30_1920 VDD VSS sg13g2_FILL8
XSTDFILL30_1928 VDD VSS sg13g2_FILL8
XSTDFILL30_1936 VDD VSS sg13g2_FILL8
XSTDFILL30_1944 VDD VSS sg13g2_FILL8
XSTDFILL30_1952 VDD VSS sg13g2_FILL8
XSTDFILL30_1960 VDD VSS sg13g2_FILL8
XSTDFILL30_1968 VDD VSS sg13g2_FILL8
XSTDFILL30_1976 VDD VSS sg13g2_FILL8
XSTDFILL30_1984 VDD VSS sg13g2_FILL8
XSTDFILL30_1992 VDD VSS sg13g2_FILL8
XSTDFILL30_2000 VDD VSS sg13g2_FILL8
XSTDFILL30_2008 VDD VSS sg13g2_FILL8
XSTDFILL30_2016 VDD VSS sg13g2_FILL8
XSTDFILL30_2024 VDD VSS sg13g2_FILL8
XSTDFILL30_2032 VDD VSS sg13g2_FILL8
XSTDFILL30_2040 VDD VSS sg13g2_FILL8
XSTDFILL30_2048 VDD VSS sg13g2_FILL8
XSTDFILL30_2056 VDD VSS sg13g2_FILL8
XSTDFILL30_2064 VDD VSS sg13g2_FILL8
XSTDFILL30_2072 VDD VSS sg13g2_FILL8
XSTDFILL30_2080 VDD VSS sg13g2_FILL8
XSTDFILL30_2088 VDD VSS sg13g2_FILL8
XSTDFILL30_2096 VDD VSS sg13g2_FILL8
XSTDFILL30_2104 VDD VSS sg13g2_FILL8
XSTDFILL30_2112 VDD VSS sg13g2_FILL8
XSTDFILL30_2120 VDD VSS sg13g2_FILL8
XSTDFILL30_2128 VDD VSS sg13g2_FILL8
XSTDFILL30_2136 VDD VSS sg13g2_FILL8
XSTDFILL30_2144 VDD VSS sg13g2_FILL8
XSTDFILL30_2152 VDD VSS sg13g2_FILL8
XSTDFILL30_2160 VDD VSS sg13g2_FILL8
XSTDFILL30_2168 VDD VSS sg13g2_FILL4
XSTDFILL31_0 VDD VSS sg13g2_FILL8
XSTDFILL31_8 VDD VSS sg13g2_FILL8
XSTDFILL31_16 VDD VSS sg13g2_FILL8
XSTDFILL31_24 VDD VSS sg13g2_FILL8
XSTDFILL31_32 VDD VSS sg13g2_FILL8
XSTDFILL31_40 VDD VSS sg13g2_FILL8
XSTDFILL31_48 VDD VSS sg13g2_FILL8
XSTDFILL31_56 VDD VSS sg13g2_FILL8
XSTDFILL31_64 VDD VSS sg13g2_FILL8
XSTDFILL31_72 VDD VSS sg13g2_FILL8
XSTDFILL31_80 VDD VSS sg13g2_FILL8
XSTDFILL31_88 VDD VSS sg13g2_FILL8
XSTDFILL31_96 VDD VSS sg13g2_FILL8
XSTDFILL31_104 VDD VSS sg13g2_FILL1
XSTDFILL31_1880 VDD VSS sg13g2_FILL8
XSTDFILL31_1888 VDD VSS sg13g2_FILL8
XSTDFILL31_1896 VDD VSS sg13g2_FILL8
XSTDFILL31_1904 VDD VSS sg13g2_FILL8
XSTDFILL31_1912 VDD VSS sg13g2_FILL8
XSTDFILL31_1920 VDD VSS sg13g2_FILL8
XSTDFILL31_1928 VDD VSS sg13g2_FILL8
XSTDFILL31_1936 VDD VSS sg13g2_FILL8
XSTDFILL31_1944 VDD VSS sg13g2_FILL8
XSTDFILL31_1952 VDD VSS sg13g2_FILL8
XSTDFILL31_1960 VDD VSS sg13g2_FILL8
XSTDFILL31_1968 VDD VSS sg13g2_FILL8
XSTDFILL31_1976 VDD VSS sg13g2_FILL8
XSTDFILL31_1984 VDD VSS sg13g2_FILL8
XSTDFILL31_1992 VDD VSS sg13g2_FILL8
XSTDFILL31_2000 VDD VSS sg13g2_FILL8
XSTDFILL31_2008 VDD VSS sg13g2_FILL8
XSTDFILL31_2016 VDD VSS sg13g2_FILL8
XSTDFILL31_2024 VDD VSS sg13g2_FILL8
XSTDFILL31_2032 VDD VSS sg13g2_FILL8
XSTDFILL31_2040 VDD VSS sg13g2_FILL8
XSTDFILL31_2048 VDD VSS sg13g2_FILL8
XSTDFILL31_2056 VDD VSS sg13g2_FILL8
XSTDFILL31_2064 VDD VSS sg13g2_FILL8
XSTDFILL31_2072 VDD VSS sg13g2_FILL8
XSTDFILL31_2080 VDD VSS sg13g2_FILL8
XSTDFILL31_2088 VDD VSS sg13g2_FILL8
XSTDFILL31_2096 VDD VSS sg13g2_FILL8
XSTDFILL31_2104 VDD VSS sg13g2_FILL8
XSTDFILL31_2112 VDD VSS sg13g2_FILL8
XSTDFILL31_2120 VDD VSS sg13g2_FILL8
XSTDFILL31_2128 VDD VSS sg13g2_FILL8
XSTDFILL31_2136 VDD VSS sg13g2_FILL8
XSTDFILL31_2144 VDD VSS sg13g2_FILL8
XSTDFILL31_2152 VDD VSS sg13g2_FILL8
XSTDFILL31_2160 VDD VSS sg13g2_FILL8
XSTDFILL31_2168 VDD VSS sg13g2_FILL4
XSTDFILL32_0 VDD VSS sg13g2_FILL8
XSTDFILL32_8 VDD VSS sg13g2_FILL8
XSTDFILL32_16 VDD VSS sg13g2_FILL8
XSTDFILL32_24 VDD VSS sg13g2_FILL8
XSTDFILL32_32 VDD VSS sg13g2_FILL8
XSTDFILL32_40 VDD VSS sg13g2_FILL8
XSTDFILL32_48 VDD VSS sg13g2_FILL8
XSTDFILL32_56 VDD VSS sg13g2_FILL8
XSTDFILL32_64 VDD VSS sg13g2_FILL8
XSTDFILL32_72 VDD VSS sg13g2_FILL8
XSTDFILL32_80 VDD VSS sg13g2_FILL8
XSTDFILL32_88 VDD VSS sg13g2_FILL8
XSTDFILL32_96 VDD VSS sg13g2_FILL8
XSTDFILL32_104 VDD VSS sg13g2_FILL1
XSTDFILL32_1880 VDD VSS sg13g2_FILL8
XSTDFILL32_1888 VDD VSS sg13g2_FILL8
XSTDFILL32_1896 VDD VSS sg13g2_FILL8
XSTDFILL32_1904 VDD VSS sg13g2_FILL8
XSTDFILL32_1912 VDD VSS sg13g2_FILL8
XSTDFILL32_1920 VDD VSS sg13g2_FILL8
XSTDFILL32_1928 VDD VSS sg13g2_FILL8
XSTDFILL32_1936 VDD VSS sg13g2_FILL8
XSTDFILL32_1944 VDD VSS sg13g2_FILL8
XSTDFILL32_1952 VDD VSS sg13g2_FILL8
XSTDFILL32_1960 VDD VSS sg13g2_FILL8
XSTDFILL32_1968 VDD VSS sg13g2_FILL8
XSTDFILL32_1976 VDD VSS sg13g2_FILL8
XSTDFILL32_1984 VDD VSS sg13g2_FILL8
XSTDFILL32_1992 VDD VSS sg13g2_FILL8
XSTDFILL32_2000 VDD VSS sg13g2_FILL8
XSTDFILL32_2008 VDD VSS sg13g2_FILL8
XSTDFILL32_2016 VDD VSS sg13g2_FILL8
XSTDFILL32_2024 VDD VSS sg13g2_FILL8
XSTDFILL32_2032 VDD VSS sg13g2_FILL8
XSTDFILL32_2040 VDD VSS sg13g2_FILL8
XSTDFILL32_2048 VDD VSS sg13g2_FILL8
XSTDFILL32_2056 VDD VSS sg13g2_FILL8
XSTDFILL32_2064 VDD VSS sg13g2_FILL8
XSTDFILL32_2072 VDD VSS sg13g2_FILL8
XSTDFILL32_2080 VDD VSS sg13g2_FILL8
XSTDFILL32_2088 VDD VSS sg13g2_FILL8
XSTDFILL32_2096 VDD VSS sg13g2_FILL8
XSTDFILL32_2104 VDD VSS sg13g2_FILL8
XSTDFILL32_2112 VDD VSS sg13g2_FILL8
XSTDFILL32_2120 VDD VSS sg13g2_FILL8
XSTDFILL32_2128 VDD VSS sg13g2_FILL8
XSTDFILL32_2136 VDD VSS sg13g2_FILL8
XSTDFILL32_2144 VDD VSS sg13g2_FILL8
XSTDFILL32_2152 VDD VSS sg13g2_FILL8
XSTDFILL32_2160 VDD VSS sg13g2_FILL8
XSTDFILL32_2168 VDD VSS sg13g2_FILL4
XSTDFILL33_0 VDD VSS sg13g2_FILL8
XSTDFILL33_8 VDD VSS sg13g2_FILL8
XSTDFILL33_16 VDD VSS sg13g2_FILL8
XSTDFILL33_24 VDD VSS sg13g2_FILL8
XSTDFILL33_32 VDD VSS sg13g2_FILL8
XSTDFILL33_40 VDD VSS sg13g2_FILL8
XSTDFILL33_48 VDD VSS sg13g2_FILL8
XSTDFILL33_56 VDD VSS sg13g2_FILL8
XSTDFILL33_64 VDD VSS sg13g2_FILL8
XSTDFILL33_72 VDD VSS sg13g2_FILL8
XSTDFILL33_80 VDD VSS sg13g2_FILL8
XSTDFILL33_88 VDD VSS sg13g2_FILL8
XSTDFILL33_96 VDD VSS sg13g2_FILL8
XSTDFILL33_104 VDD VSS sg13g2_FILL1
XSTDFILL33_1880 VDD VSS sg13g2_FILL8
XSTDFILL33_1888 VDD VSS sg13g2_FILL8
XSTDFILL33_1896 VDD VSS sg13g2_FILL8
XSTDFILL33_1904 VDD VSS sg13g2_FILL8
XSTDFILL33_1912 VDD VSS sg13g2_FILL8
XSTDFILL33_1920 VDD VSS sg13g2_FILL8
XSTDFILL33_1928 VDD VSS sg13g2_FILL8
XSTDFILL33_1936 VDD VSS sg13g2_FILL8
XSTDFILL33_1944 VDD VSS sg13g2_FILL8
XSTDFILL33_1952 VDD VSS sg13g2_FILL8
XSTDFILL33_1960 VDD VSS sg13g2_FILL8
XSTDFILL33_1968 VDD VSS sg13g2_FILL8
XSTDFILL33_1976 VDD VSS sg13g2_FILL8
XSTDFILL33_1984 VDD VSS sg13g2_FILL8
XSTDFILL33_1992 VDD VSS sg13g2_FILL8
XSTDFILL33_2000 VDD VSS sg13g2_FILL8
XSTDFILL33_2008 VDD VSS sg13g2_FILL8
XSTDFILL33_2016 VDD VSS sg13g2_FILL8
XSTDFILL33_2024 VDD VSS sg13g2_FILL8
XSTDFILL33_2032 VDD VSS sg13g2_FILL8
XSTDFILL33_2040 VDD VSS sg13g2_FILL8
XSTDFILL33_2048 VDD VSS sg13g2_FILL8
XSTDFILL33_2056 VDD VSS sg13g2_FILL8
XSTDFILL33_2064 VDD VSS sg13g2_FILL8
XSTDFILL33_2072 VDD VSS sg13g2_FILL8
XSTDFILL33_2080 VDD VSS sg13g2_FILL8
XSTDFILL33_2088 VDD VSS sg13g2_FILL8
XSTDFILL33_2096 VDD VSS sg13g2_FILL8
XSTDFILL33_2104 VDD VSS sg13g2_FILL8
XSTDFILL33_2112 VDD VSS sg13g2_FILL8
XSTDFILL33_2120 VDD VSS sg13g2_FILL8
XSTDFILL33_2128 VDD VSS sg13g2_FILL8
XSTDFILL33_2136 VDD VSS sg13g2_FILL8
XSTDFILL33_2144 VDD VSS sg13g2_FILL8
XSTDFILL33_2152 VDD VSS sg13g2_FILL8
XSTDFILL33_2160 VDD VSS sg13g2_FILL8
XSTDFILL33_2168 VDD VSS sg13g2_FILL4
XSTDFILL34_0 VDD VSS sg13g2_FILL8
XSTDFILL34_8 VDD VSS sg13g2_FILL8
XSTDFILL34_16 VDD VSS sg13g2_FILL8
XSTDFILL34_24 VDD VSS sg13g2_FILL8
XSTDFILL34_32 VDD VSS sg13g2_FILL8
XSTDFILL34_40 VDD VSS sg13g2_FILL8
XSTDFILL34_48 VDD VSS sg13g2_FILL8
XSTDFILL34_56 VDD VSS sg13g2_FILL8
XSTDFILL34_64 VDD VSS sg13g2_FILL8
XSTDFILL34_72 VDD VSS sg13g2_FILL8
XSTDFILL34_80 VDD VSS sg13g2_FILL8
XSTDFILL34_88 VDD VSS sg13g2_FILL8
XSTDFILL34_96 VDD VSS sg13g2_FILL8
XSTDFILL34_104 VDD VSS sg13g2_FILL1
XSTDFILL34_1880 VDD VSS sg13g2_FILL8
XSTDFILL34_1888 VDD VSS sg13g2_FILL8
XSTDFILL34_1896 VDD VSS sg13g2_FILL8
XSTDFILL34_1904 VDD VSS sg13g2_FILL8
XSTDFILL34_1912 VDD VSS sg13g2_FILL8
XSTDFILL34_1920 VDD VSS sg13g2_FILL8
XSTDFILL34_1928 VDD VSS sg13g2_FILL8
XSTDFILL34_1936 VDD VSS sg13g2_FILL8
XSTDFILL34_1944 VDD VSS sg13g2_FILL8
XSTDFILL34_1952 VDD VSS sg13g2_FILL8
XSTDFILL34_1960 VDD VSS sg13g2_FILL8
XSTDFILL34_1968 VDD VSS sg13g2_FILL8
XSTDFILL34_1976 VDD VSS sg13g2_FILL8
XSTDFILL34_1984 VDD VSS sg13g2_FILL8
XSTDFILL34_1992 VDD VSS sg13g2_FILL8
XSTDFILL34_2000 VDD VSS sg13g2_FILL8
XSTDFILL34_2008 VDD VSS sg13g2_FILL8
XSTDFILL34_2016 VDD VSS sg13g2_FILL8
XSTDFILL34_2024 VDD VSS sg13g2_FILL8
XSTDFILL34_2032 VDD VSS sg13g2_FILL8
XSTDFILL34_2040 VDD VSS sg13g2_FILL8
XSTDFILL34_2048 VDD VSS sg13g2_FILL8
XSTDFILL34_2056 VDD VSS sg13g2_FILL8
XSTDFILL34_2064 VDD VSS sg13g2_FILL8
XSTDFILL34_2072 VDD VSS sg13g2_FILL8
XSTDFILL34_2080 VDD VSS sg13g2_FILL8
XSTDFILL34_2088 VDD VSS sg13g2_FILL8
XSTDFILL34_2096 VDD VSS sg13g2_FILL8
XSTDFILL34_2104 VDD VSS sg13g2_FILL8
XSTDFILL34_2112 VDD VSS sg13g2_FILL8
XSTDFILL34_2120 VDD VSS sg13g2_FILL8
XSTDFILL34_2128 VDD VSS sg13g2_FILL8
XSTDFILL34_2136 VDD VSS sg13g2_FILL8
XSTDFILL34_2144 VDD VSS sg13g2_FILL8
XSTDFILL34_2152 VDD VSS sg13g2_FILL8
XSTDFILL34_2160 VDD VSS sg13g2_FILL8
XSTDFILL34_2168 VDD VSS sg13g2_FILL4
XSTDFILL35_0 VDD VSS sg13g2_FILL8
XSTDFILL35_8 VDD VSS sg13g2_FILL8
XSTDFILL35_16 VDD VSS sg13g2_FILL8
XSTDFILL35_24 VDD VSS sg13g2_FILL8
XSTDFILL35_32 VDD VSS sg13g2_FILL8
XSTDFILL35_40 VDD VSS sg13g2_FILL8
XSTDFILL35_48 VDD VSS sg13g2_FILL8
XSTDFILL35_56 VDD VSS sg13g2_FILL8
XSTDFILL35_64 VDD VSS sg13g2_FILL8
XSTDFILL35_72 VDD VSS sg13g2_FILL8
XSTDFILL35_80 VDD VSS sg13g2_FILL8
XSTDFILL35_88 VDD VSS sg13g2_FILL8
XSTDFILL35_96 VDD VSS sg13g2_FILL8
XSTDFILL35_104 VDD VSS sg13g2_FILL1
XSTDFILL35_1880 VDD VSS sg13g2_FILL8
XSTDFILL35_1888 VDD VSS sg13g2_FILL8
XSTDFILL35_1896 VDD VSS sg13g2_FILL8
XSTDFILL35_1904 VDD VSS sg13g2_FILL8
XSTDFILL35_1912 VDD VSS sg13g2_FILL8
XSTDFILL35_1920 VDD VSS sg13g2_FILL8
XSTDFILL35_1928 VDD VSS sg13g2_FILL8
XSTDFILL35_1936 VDD VSS sg13g2_FILL8
XSTDFILL35_1944 VDD VSS sg13g2_FILL8
XSTDFILL35_1952 VDD VSS sg13g2_FILL8
XSTDFILL35_1960 VDD VSS sg13g2_FILL8
XSTDFILL35_1968 VDD VSS sg13g2_FILL8
XSTDFILL35_1976 VDD VSS sg13g2_FILL8
XSTDFILL35_1984 VDD VSS sg13g2_FILL8
XSTDFILL35_1992 VDD VSS sg13g2_FILL8
XSTDFILL35_2000 VDD VSS sg13g2_FILL8
XSTDFILL35_2008 VDD VSS sg13g2_FILL8
XSTDFILL35_2016 VDD VSS sg13g2_FILL8
XSTDFILL35_2024 VDD VSS sg13g2_FILL8
XSTDFILL35_2032 VDD VSS sg13g2_FILL8
XSTDFILL35_2040 VDD VSS sg13g2_FILL8
XSTDFILL35_2048 VDD VSS sg13g2_FILL8
XSTDFILL35_2056 VDD VSS sg13g2_FILL8
XSTDFILL35_2064 VDD VSS sg13g2_FILL8
XSTDFILL35_2072 VDD VSS sg13g2_FILL8
XSTDFILL35_2080 VDD VSS sg13g2_FILL8
XSTDFILL35_2088 VDD VSS sg13g2_FILL8
XSTDFILL35_2096 VDD VSS sg13g2_FILL8
XSTDFILL35_2104 VDD VSS sg13g2_FILL8
XSTDFILL35_2112 VDD VSS sg13g2_FILL8
XSTDFILL35_2120 VDD VSS sg13g2_FILL8
XSTDFILL35_2128 VDD VSS sg13g2_FILL8
XSTDFILL35_2136 VDD VSS sg13g2_FILL8
XSTDFILL35_2144 VDD VSS sg13g2_FILL8
XSTDFILL35_2152 VDD VSS sg13g2_FILL8
XSTDFILL35_2160 VDD VSS sg13g2_FILL8
XSTDFILL35_2168 VDD VSS sg13g2_FILL4
XSTDFILL36_0 VDD VSS sg13g2_FILL8
XSTDFILL36_8 VDD VSS sg13g2_FILL8
XSTDFILL36_16 VDD VSS sg13g2_FILL8
XSTDFILL36_24 VDD VSS sg13g2_FILL8
XSTDFILL36_32 VDD VSS sg13g2_FILL8
XSTDFILL36_40 VDD VSS sg13g2_FILL8
XSTDFILL36_48 VDD VSS sg13g2_FILL8
XSTDFILL36_56 VDD VSS sg13g2_FILL8
XSTDFILL36_64 VDD VSS sg13g2_FILL8
XSTDFILL36_72 VDD VSS sg13g2_FILL8
XSTDFILL36_80 VDD VSS sg13g2_FILL8
XSTDFILL36_88 VDD VSS sg13g2_FILL8
XSTDFILL36_96 VDD VSS sg13g2_FILL8
XSTDFILL36_104 VDD VSS sg13g2_FILL1
XSTDFILL36_1880 VDD VSS sg13g2_FILL8
XSTDFILL36_1888 VDD VSS sg13g2_FILL8
XSTDFILL36_1896 VDD VSS sg13g2_FILL8
XSTDFILL36_1904 VDD VSS sg13g2_FILL8
XSTDFILL36_1912 VDD VSS sg13g2_FILL8
XSTDFILL36_1920 VDD VSS sg13g2_FILL8
XSTDFILL36_1928 VDD VSS sg13g2_FILL8
XSTDFILL36_1936 VDD VSS sg13g2_FILL8
XSTDFILL36_1944 VDD VSS sg13g2_FILL8
XSTDFILL36_1952 VDD VSS sg13g2_FILL8
XSTDFILL36_1960 VDD VSS sg13g2_FILL8
XSTDFILL36_1968 VDD VSS sg13g2_FILL8
XSTDFILL36_1976 VDD VSS sg13g2_FILL8
XSTDFILL36_1984 VDD VSS sg13g2_FILL8
XSTDFILL36_1992 VDD VSS sg13g2_FILL8
XSTDFILL36_2000 VDD VSS sg13g2_FILL8
XSTDFILL36_2008 VDD VSS sg13g2_FILL8
XSTDFILL36_2016 VDD VSS sg13g2_FILL8
XSTDFILL36_2024 VDD VSS sg13g2_FILL8
XSTDFILL36_2032 VDD VSS sg13g2_FILL8
XSTDFILL36_2040 VDD VSS sg13g2_FILL8
XSTDFILL36_2048 VDD VSS sg13g2_FILL8
XSTDFILL36_2056 VDD VSS sg13g2_FILL8
XSTDFILL36_2064 VDD VSS sg13g2_FILL8
XSTDFILL36_2072 VDD VSS sg13g2_FILL8
XSTDFILL36_2080 VDD VSS sg13g2_FILL8
XSTDFILL36_2088 VDD VSS sg13g2_FILL8
XSTDFILL36_2096 VDD VSS sg13g2_FILL8
XSTDFILL36_2104 VDD VSS sg13g2_FILL8
XSTDFILL36_2112 VDD VSS sg13g2_FILL8
XSTDFILL36_2120 VDD VSS sg13g2_FILL8
XSTDFILL36_2128 VDD VSS sg13g2_FILL8
XSTDFILL36_2136 VDD VSS sg13g2_FILL8
XSTDFILL36_2144 VDD VSS sg13g2_FILL8
XSTDFILL36_2152 VDD VSS sg13g2_FILL8
XSTDFILL36_2160 VDD VSS sg13g2_FILL8
XSTDFILL36_2168 VDD VSS sg13g2_FILL4
XSTDFILL37_0 VDD VSS sg13g2_FILL8
XSTDFILL37_8 VDD VSS sg13g2_FILL8
XSTDFILL37_16 VDD VSS sg13g2_FILL8
XSTDFILL37_24 VDD VSS sg13g2_FILL8
XSTDFILL37_32 VDD VSS sg13g2_FILL8
XSTDFILL37_40 VDD VSS sg13g2_FILL8
XSTDFILL37_48 VDD VSS sg13g2_FILL8
XSTDFILL37_56 VDD VSS sg13g2_FILL8
XSTDFILL37_64 VDD VSS sg13g2_FILL8
XSTDFILL37_72 VDD VSS sg13g2_FILL8
XSTDFILL37_80 VDD VSS sg13g2_FILL8
XSTDFILL37_88 VDD VSS sg13g2_FILL8
XSTDFILL37_96 VDD VSS sg13g2_FILL8
XSTDFILL37_104 VDD VSS sg13g2_FILL1
XSTDFILL37_1880 VDD VSS sg13g2_FILL8
XSTDFILL37_1888 VDD VSS sg13g2_FILL8
XSTDFILL37_1896 VDD VSS sg13g2_FILL8
XSTDFILL37_1904 VDD VSS sg13g2_FILL8
XSTDFILL37_1912 VDD VSS sg13g2_FILL8
XSTDFILL37_1920 VDD VSS sg13g2_FILL8
XSTDFILL37_1928 VDD VSS sg13g2_FILL8
XSTDFILL37_1936 VDD VSS sg13g2_FILL8
XSTDFILL37_1944 VDD VSS sg13g2_FILL8
XSTDFILL37_1952 VDD VSS sg13g2_FILL8
XSTDFILL37_1960 VDD VSS sg13g2_FILL8
XSTDFILL37_1968 VDD VSS sg13g2_FILL8
XSTDFILL37_1976 VDD VSS sg13g2_FILL8
XSTDFILL37_1984 VDD VSS sg13g2_FILL8
XSTDFILL37_1992 VDD VSS sg13g2_FILL8
XSTDFILL37_2000 VDD VSS sg13g2_FILL8
XSTDFILL37_2008 VDD VSS sg13g2_FILL8
XSTDFILL37_2016 VDD VSS sg13g2_FILL8
XSTDFILL37_2024 VDD VSS sg13g2_FILL8
XSTDFILL37_2032 VDD VSS sg13g2_FILL8
XSTDFILL37_2040 VDD VSS sg13g2_FILL8
XSTDFILL37_2048 VDD VSS sg13g2_FILL8
XSTDFILL37_2056 VDD VSS sg13g2_FILL8
XSTDFILL37_2064 VDD VSS sg13g2_FILL8
XSTDFILL37_2072 VDD VSS sg13g2_FILL8
XSTDFILL37_2080 VDD VSS sg13g2_FILL8
XSTDFILL37_2088 VDD VSS sg13g2_FILL8
XSTDFILL37_2096 VDD VSS sg13g2_FILL8
XSTDFILL37_2104 VDD VSS sg13g2_FILL8
XSTDFILL37_2112 VDD VSS sg13g2_FILL8
XSTDFILL37_2120 VDD VSS sg13g2_FILL8
XSTDFILL37_2128 VDD VSS sg13g2_FILL8
XSTDFILL37_2136 VDD VSS sg13g2_FILL8
XSTDFILL37_2144 VDD VSS sg13g2_FILL8
XSTDFILL37_2152 VDD VSS sg13g2_FILL8
XSTDFILL37_2160 VDD VSS sg13g2_FILL8
XSTDFILL37_2168 VDD VSS sg13g2_FILL4
XSTDFILL38_0 VDD VSS sg13g2_FILL8
XSTDFILL38_8 VDD VSS sg13g2_FILL8
XSTDFILL38_16 VDD VSS sg13g2_FILL8
XSTDFILL38_24 VDD VSS sg13g2_FILL8
XSTDFILL38_32 VDD VSS sg13g2_FILL8
XSTDFILL38_40 VDD VSS sg13g2_FILL8
XSTDFILL38_48 VDD VSS sg13g2_FILL8
XSTDFILL38_56 VDD VSS sg13g2_FILL8
XSTDFILL38_64 VDD VSS sg13g2_FILL8
XSTDFILL38_72 VDD VSS sg13g2_FILL8
XSTDFILL38_80 VDD VSS sg13g2_FILL8
XSTDFILL38_88 VDD VSS sg13g2_FILL8
XSTDFILL38_96 VDD VSS sg13g2_FILL8
XSTDFILL38_104 VDD VSS sg13g2_FILL1
XSTDFILL38_1880 VDD VSS sg13g2_FILL8
XSTDFILL38_1888 VDD VSS sg13g2_FILL8
XSTDFILL38_1896 VDD VSS sg13g2_FILL8
XSTDFILL38_1904 VDD VSS sg13g2_FILL8
XSTDFILL38_1912 VDD VSS sg13g2_FILL8
XSTDFILL38_1920 VDD VSS sg13g2_FILL8
XSTDFILL38_1928 VDD VSS sg13g2_FILL8
XSTDFILL38_1936 VDD VSS sg13g2_FILL8
XSTDFILL38_1944 VDD VSS sg13g2_FILL8
XSTDFILL38_1952 VDD VSS sg13g2_FILL8
XSTDFILL38_1960 VDD VSS sg13g2_FILL8
XSTDFILL38_1968 VDD VSS sg13g2_FILL8
XSTDFILL38_1976 VDD VSS sg13g2_FILL8
XSTDFILL38_1984 VDD VSS sg13g2_FILL8
XSTDFILL38_1992 VDD VSS sg13g2_FILL8
XSTDFILL38_2000 VDD VSS sg13g2_FILL8
XSTDFILL38_2008 VDD VSS sg13g2_FILL8
XSTDFILL38_2016 VDD VSS sg13g2_FILL8
XSTDFILL38_2024 VDD VSS sg13g2_FILL8
XSTDFILL38_2032 VDD VSS sg13g2_FILL8
XSTDFILL38_2040 VDD VSS sg13g2_FILL8
XSTDFILL38_2048 VDD VSS sg13g2_FILL8
XSTDFILL38_2056 VDD VSS sg13g2_FILL8
XSTDFILL38_2064 VDD VSS sg13g2_FILL8
XSTDFILL38_2072 VDD VSS sg13g2_FILL8
XSTDFILL38_2080 VDD VSS sg13g2_FILL8
XSTDFILL38_2088 VDD VSS sg13g2_FILL8
XSTDFILL38_2096 VDD VSS sg13g2_FILL8
XSTDFILL38_2104 VDD VSS sg13g2_FILL8
XSTDFILL38_2112 VDD VSS sg13g2_FILL8
XSTDFILL38_2120 VDD VSS sg13g2_FILL8
XSTDFILL38_2128 VDD VSS sg13g2_FILL8
XSTDFILL38_2136 VDD VSS sg13g2_FILL8
XSTDFILL38_2144 VDD VSS sg13g2_FILL8
XSTDFILL38_2152 VDD VSS sg13g2_FILL8
XSTDFILL38_2160 VDD VSS sg13g2_FILL8
XSTDFILL38_2168 VDD VSS sg13g2_FILL4
XSTDFILL39_0 VDD VSS sg13g2_FILL8
XSTDFILL39_8 VDD VSS sg13g2_FILL8
XSTDFILL39_16 VDD VSS sg13g2_FILL8
XSTDFILL39_24 VDD VSS sg13g2_FILL8
XSTDFILL39_32 VDD VSS sg13g2_FILL8
XSTDFILL39_40 VDD VSS sg13g2_FILL8
XSTDFILL39_48 VDD VSS sg13g2_FILL8
XSTDFILL39_56 VDD VSS sg13g2_FILL8
XSTDFILL39_64 VDD VSS sg13g2_FILL8
XSTDFILL39_72 VDD VSS sg13g2_FILL8
XSTDFILL39_80 VDD VSS sg13g2_FILL8
XSTDFILL39_88 VDD VSS sg13g2_FILL8
XSTDFILL39_96 VDD VSS sg13g2_FILL8
XSTDFILL39_104 VDD VSS sg13g2_FILL1
XSTDFILL39_1880 VDD VSS sg13g2_FILL8
XSTDFILL39_1888 VDD VSS sg13g2_FILL8
XSTDFILL39_1896 VDD VSS sg13g2_FILL8
XSTDFILL39_1904 VDD VSS sg13g2_FILL8
XSTDFILL39_1912 VDD VSS sg13g2_FILL8
XSTDFILL39_1920 VDD VSS sg13g2_FILL8
XSTDFILL39_1928 VDD VSS sg13g2_FILL8
XSTDFILL39_1936 VDD VSS sg13g2_FILL8
XSTDFILL39_1944 VDD VSS sg13g2_FILL8
XSTDFILL39_1952 VDD VSS sg13g2_FILL8
XSTDFILL39_1960 VDD VSS sg13g2_FILL8
XSTDFILL39_1968 VDD VSS sg13g2_FILL8
XSTDFILL39_1976 VDD VSS sg13g2_FILL8
XSTDFILL39_1984 VDD VSS sg13g2_FILL8
XSTDFILL39_1992 VDD VSS sg13g2_FILL8
XSTDFILL39_2000 VDD VSS sg13g2_FILL8
XSTDFILL39_2008 VDD VSS sg13g2_FILL8
XSTDFILL39_2016 VDD VSS sg13g2_FILL8
XSTDFILL39_2024 VDD VSS sg13g2_FILL8
XSTDFILL39_2032 VDD VSS sg13g2_FILL8
XSTDFILL39_2040 VDD VSS sg13g2_FILL8
XSTDFILL39_2048 VDD VSS sg13g2_FILL8
XSTDFILL39_2056 VDD VSS sg13g2_FILL8
XSTDFILL39_2064 VDD VSS sg13g2_FILL8
XSTDFILL39_2072 VDD VSS sg13g2_FILL8
XSTDFILL39_2080 VDD VSS sg13g2_FILL8
XSTDFILL39_2088 VDD VSS sg13g2_FILL8
XSTDFILL39_2096 VDD VSS sg13g2_FILL8
XSTDFILL39_2104 VDD VSS sg13g2_FILL8
XSTDFILL39_2112 VDD VSS sg13g2_FILL8
XSTDFILL39_2120 VDD VSS sg13g2_FILL8
XSTDFILL39_2128 VDD VSS sg13g2_FILL8
XSTDFILL39_2136 VDD VSS sg13g2_FILL8
XSTDFILL39_2144 VDD VSS sg13g2_FILL8
XSTDFILL39_2152 VDD VSS sg13g2_FILL8
XSTDFILL39_2160 VDD VSS sg13g2_FILL8
XSTDFILL39_2168 VDD VSS sg13g2_FILL4
XSTDFILL40_0 VDD VSS sg13g2_FILL8
XSTDFILL40_8 VDD VSS sg13g2_FILL8
XSTDFILL40_16 VDD VSS sg13g2_FILL8
XSTDFILL40_24 VDD VSS sg13g2_FILL8
XSTDFILL40_32 VDD VSS sg13g2_FILL8
XSTDFILL40_40 VDD VSS sg13g2_FILL8
XSTDFILL40_48 VDD VSS sg13g2_FILL8
XSTDFILL40_56 VDD VSS sg13g2_FILL8
XSTDFILL40_64 VDD VSS sg13g2_FILL8
XSTDFILL40_72 VDD VSS sg13g2_FILL8
XSTDFILL40_80 VDD VSS sg13g2_FILL8
XSTDFILL40_88 VDD VSS sg13g2_FILL8
XSTDFILL40_96 VDD VSS sg13g2_FILL8
XSTDFILL40_104 VDD VSS sg13g2_FILL1
XSTDFILL40_1880 VDD VSS sg13g2_FILL8
XSTDFILL40_1888 VDD VSS sg13g2_FILL8
XSTDFILL40_1896 VDD VSS sg13g2_FILL8
XSTDFILL40_1904 VDD VSS sg13g2_FILL8
XSTDFILL40_1912 VDD VSS sg13g2_FILL8
XSTDFILL40_1920 VDD VSS sg13g2_FILL8
XSTDFILL40_1928 VDD VSS sg13g2_FILL8
XSTDFILL40_1936 VDD VSS sg13g2_FILL8
XSTDFILL40_1944 VDD VSS sg13g2_FILL8
XSTDFILL40_1952 VDD VSS sg13g2_FILL8
XSTDFILL40_1960 VDD VSS sg13g2_FILL8
XSTDFILL40_1968 VDD VSS sg13g2_FILL8
XSTDFILL40_1976 VDD VSS sg13g2_FILL8
XSTDFILL40_1984 VDD VSS sg13g2_FILL8
XSTDFILL40_1992 VDD VSS sg13g2_FILL8
XSTDFILL40_2000 VDD VSS sg13g2_FILL8
XSTDFILL40_2008 VDD VSS sg13g2_FILL8
XSTDFILL40_2016 VDD VSS sg13g2_FILL8
XSTDFILL40_2024 VDD VSS sg13g2_FILL8
XSTDFILL40_2032 VDD VSS sg13g2_FILL8
XSTDFILL40_2040 VDD VSS sg13g2_FILL8
XSTDFILL40_2048 VDD VSS sg13g2_FILL8
XSTDFILL40_2056 VDD VSS sg13g2_FILL8
XSTDFILL40_2064 VDD VSS sg13g2_FILL8
XSTDFILL40_2072 VDD VSS sg13g2_FILL8
XSTDFILL40_2080 VDD VSS sg13g2_FILL8
XSTDFILL40_2088 VDD VSS sg13g2_FILL8
XSTDFILL40_2096 VDD VSS sg13g2_FILL8
XSTDFILL40_2104 VDD VSS sg13g2_FILL8
XSTDFILL40_2112 VDD VSS sg13g2_FILL8
XSTDFILL40_2120 VDD VSS sg13g2_FILL8
XSTDFILL40_2128 VDD VSS sg13g2_FILL8
XSTDFILL40_2136 VDD VSS sg13g2_FILL8
XSTDFILL40_2144 VDD VSS sg13g2_FILL8
XSTDFILL40_2152 VDD VSS sg13g2_FILL8
XSTDFILL40_2160 VDD VSS sg13g2_FILL8
XSTDFILL40_2168 VDD VSS sg13g2_FILL4
XSTDFILL41_0 VDD VSS sg13g2_FILL8
XSTDFILL41_8 VDD VSS sg13g2_FILL8
XSTDFILL41_16 VDD VSS sg13g2_FILL8
XSTDFILL41_24 VDD VSS sg13g2_FILL8
XSTDFILL41_32 VDD VSS sg13g2_FILL8
XSTDFILL41_40 VDD VSS sg13g2_FILL8
XSTDFILL41_48 VDD VSS sg13g2_FILL8
XSTDFILL41_56 VDD VSS sg13g2_FILL8
XSTDFILL41_64 VDD VSS sg13g2_FILL8
XSTDFILL41_72 VDD VSS sg13g2_FILL8
XSTDFILL41_80 VDD VSS sg13g2_FILL8
XSTDFILL41_88 VDD VSS sg13g2_FILL8
XSTDFILL41_96 VDD VSS sg13g2_FILL8
XSTDFILL41_104 VDD VSS sg13g2_FILL1
XSTDFILL41_1880 VDD VSS sg13g2_FILL8
XSTDFILL41_1888 VDD VSS sg13g2_FILL8
XSTDFILL41_1896 VDD VSS sg13g2_FILL8
XSTDFILL41_1904 VDD VSS sg13g2_FILL8
XSTDFILL41_1912 VDD VSS sg13g2_FILL8
XSTDFILL41_1920 VDD VSS sg13g2_FILL8
XSTDFILL41_1928 VDD VSS sg13g2_FILL8
XSTDFILL41_1936 VDD VSS sg13g2_FILL8
XSTDFILL41_1944 VDD VSS sg13g2_FILL8
XSTDFILL41_1952 VDD VSS sg13g2_FILL8
XSTDFILL41_1960 VDD VSS sg13g2_FILL8
XSTDFILL41_1968 VDD VSS sg13g2_FILL8
XSTDFILL41_1976 VDD VSS sg13g2_FILL8
XSTDFILL41_1984 VDD VSS sg13g2_FILL8
XSTDFILL41_1992 VDD VSS sg13g2_FILL8
XSTDFILL41_2000 VDD VSS sg13g2_FILL8
XSTDFILL41_2008 VDD VSS sg13g2_FILL8
XSTDFILL41_2016 VDD VSS sg13g2_FILL8
XSTDFILL41_2024 VDD VSS sg13g2_FILL8
XSTDFILL41_2032 VDD VSS sg13g2_FILL8
XSTDFILL41_2040 VDD VSS sg13g2_FILL8
XSTDFILL41_2048 VDD VSS sg13g2_FILL8
XSTDFILL41_2056 VDD VSS sg13g2_FILL8
XSTDFILL41_2064 VDD VSS sg13g2_FILL8
XSTDFILL41_2072 VDD VSS sg13g2_FILL8
XSTDFILL41_2080 VDD VSS sg13g2_FILL8
XSTDFILL41_2088 VDD VSS sg13g2_FILL8
XSTDFILL41_2096 VDD VSS sg13g2_FILL8
XSTDFILL41_2104 VDD VSS sg13g2_FILL8
XSTDFILL41_2112 VDD VSS sg13g2_FILL8
XSTDFILL41_2120 VDD VSS sg13g2_FILL8
XSTDFILL41_2128 VDD VSS sg13g2_FILL8
XSTDFILL41_2136 VDD VSS sg13g2_FILL8
XSTDFILL41_2144 VDD VSS sg13g2_FILL8
XSTDFILL41_2152 VDD VSS sg13g2_FILL8
XSTDFILL41_2160 VDD VSS sg13g2_FILL8
XSTDFILL41_2168 VDD VSS sg13g2_FILL4
XSTDFILL42_0 VDD VSS sg13g2_FILL8
XSTDFILL42_8 VDD VSS sg13g2_FILL8
XSTDFILL42_16 VDD VSS sg13g2_FILL8
XSTDFILL42_24 VDD VSS sg13g2_FILL8
XSTDFILL42_32 VDD VSS sg13g2_FILL8
XSTDFILL42_40 VDD VSS sg13g2_FILL8
XSTDFILL42_48 VDD VSS sg13g2_FILL8
XSTDFILL42_56 VDD VSS sg13g2_FILL8
XSTDFILL42_64 VDD VSS sg13g2_FILL8
XSTDFILL42_72 VDD VSS sg13g2_FILL8
XSTDFILL42_80 VDD VSS sg13g2_FILL8
XSTDFILL42_88 VDD VSS sg13g2_FILL8
XSTDFILL42_96 VDD VSS sg13g2_FILL8
XSTDFILL42_104 VDD VSS sg13g2_FILL1
XSTDFILL42_1880 VDD VSS sg13g2_FILL8
XSTDFILL42_1888 VDD VSS sg13g2_FILL8
XSTDFILL42_1896 VDD VSS sg13g2_FILL8
XSTDFILL42_1904 VDD VSS sg13g2_FILL8
XSTDFILL42_1912 VDD VSS sg13g2_FILL8
XSTDFILL42_1920 VDD VSS sg13g2_FILL8
XSTDFILL42_1928 VDD VSS sg13g2_FILL8
XSTDFILL42_1936 VDD VSS sg13g2_FILL8
XSTDFILL42_1944 VDD VSS sg13g2_FILL8
XSTDFILL42_1952 VDD VSS sg13g2_FILL8
XSTDFILL42_1960 VDD VSS sg13g2_FILL8
XSTDFILL42_1968 VDD VSS sg13g2_FILL8
XSTDFILL42_1976 VDD VSS sg13g2_FILL8
XSTDFILL42_1984 VDD VSS sg13g2_FILL8
XSTDFILL42_1992 VDD VSS sg13g2_FILL8
XSTDFILL42_2000 VDD VSS sg13g2_FILL8
XSTDFILL42_2008 VDD VSS sg13g2_FILL8
XSTDFILL42_2016 VDD VSS sg13g2_FILL8
XSTDFILL42_2024 VDD VSS sg13g2_FILL8
XSTDFILL42_2032 VDD VSS sg13g2_FILL8
XSTDFILL42_2040 VDD VSS sg13g2_FILL8
XSTDFILL42_2048 VDD VSS sg13g2_FILL8
XSTDFILL42_2056 VDD VSS sg13g2_FILL8
XSTDFILL42_2064 VDD VSS sg13g2_FILL8
XSTDFILL42_2072 VDD VSS sg13g2_FILL8
XSTDFILL42_2080 VDD VSS sg13g2_FILL8
XSTDFILL42_2088 VDD VSS sg13g2_FILL8
XSTDFILL42_2096 VDD VSS sg13g2_FILL8
XSTDFILL42_2104 VDD VSS sg13g2_FILL8
XSTDFILL42_2112 VDD VSS sg13g2_FILL8
XSTDFILL42_2120 VDD VSS sg13g2_FILL8
XSTDFILL42_2128 VDD VSS sg13g2_FILL8
XSTDFILL42_2136 VDD VSS sg13g2_FILL8
XSTDFILL42_2144 VDD VSS sg13g2_FILL8
XSTDFILL42_2152 VDD VSS sg13g2_FILL8
XSTDFILL42_2160 VDD VSS sg13g2_FILL8
XSTDFILL42_2168 VDD VSS sg13g2_FILL4
XSTDFILL43_0 VDD VSS sg13g2_FILL8
XSTDFILL43_8 VDD VSS sg13g2_FILL8
XSTDFILL43_16 VDD VSS sg13g2_FILL8
XSTDFILL43_24 VDD VSS sg13g2_FILL8
XSTDFILL43_32 VDD VSS sg13g2_FILL8
XSTDFILL43_40 VDD VSS sg13g2_FILL8
XSTDFILL43_48 VDD VSS sg13g2_FILL8
XSTDFILL43_56 VDD VSS sg13g2_FILL8
XSTDFILL43_64 VDD VSS sg13g2_FILL8
XSTDFILL43_72 VDD VSS sg13g2_FILL8
XSTDFILL43_80 VDD VSS sg13g2_FILL8
XSTDFILL43_88 VDD VSS sg13g2_FILL8
XSTDFILL43_96 VDD VSS sg13g2_FILL8
XSTDFILL43_104 VDD VSS sg13g2_FILL1
XSTDFILL43_1880 VDD VSS sg13g2_FILL8
XSTDFILL43_1888 VDD VSS sg13g2_FILL8
XSTDFILL43_1896 VDD VSS sg13g2_FILL8
XSTDFILL43_1904 VDD VSS sg13g2_FILL8
XSTDFILL43_1912 VDD VSS sg13g2_FILL8
XSTDFILL43_1920 VDD VSS sg13g2_FILL8
XSTDFILL43_1928 VDD VSS sg13g2_FILL8
XSTDFILL43_1936 VDD VSS sg13g2_FILL8
XSTDFILL43_1944 VDD VSS sg13g2_FILL8
XSTDFILL43_1952 VDD VSS sg13g2_FILL8
XSTDFILL43_1960 VDD VSS sg13g2_FILL8
XSTDFILL43_1968 VDD VSS sg13g2_FILL8
XSTDFILL43_1976 VDD VSS sg13g2_FILL8
XSTDFILL43_1984 VDD VSS sg13g2_FILL8
XSTDFILL43_1992 VDD VSS sg13g2_FILL8
XSTDFILL43_2000 VDD VSS sg13g2_FILL8
XSTDFILL43_2008 VDD VSS sg13g2_FILL8
XSTDFILL43_2016 VDD VSS sg13g2_FILL8
XSTDFILL43_2024 VDD VSS sg13g2_FILL8
XSTDFILL43_2032 VDD VSS sg13g2_FILL8
XSTDFILL43_2040 VDD VSS sg13g2_FILL8
XSTDFILL43_2048 VDD VSS sg13g2_FILL8
XSTDFILL43_2056 VDD VSS sg13g2_FILL8
XSTDFILL43_2064 VDD VSS sg13g2_FILL8
XSTDFILL43_2072 VDD VSS sg13g2_FILL8
XSTDFILL43_2080 VDD VSS sg13g2_FILL8
XSTDFILL43_2088 VDD VSS sg13g2_FILL8
XSTDFILL43_2096 VDD VSS sg13g2_FILL8
XSTDFILL43_2104 VDD VSS sg13g2_FILL8
XSTDFILL43_2112 VDD VSS sg13g2_FILL8
XSTDFILL43_2120 VDD VSS sg13g2_FILL8
XSTDFILL43_2128 VDD VSS sg13g2_FILL8
XSTDFILL43_2136 VDD VSS sg13g2_FILL8
XSTDFILL43_2144 VDD VSS sg13g2_FILL8
XSTDFILL43_2152 VDD VSS sg13g2_FILL8
XSTDFILL43_2160 VDD VSS sg13g2_FILL8
XSTDFILL43_2168 VDD VSS sg13g2_FILL4
XSTDFILL44_0 VDD VSS sg13g2_FILL8
XSTDFILL44_8 VDD VSS sg13g2_FILL8
XSTDFILL44_16 VDD VSS sg13g2_FILL8
XSTDFILL44_24 VDD VSS sg13g2_FILL8
XSTDFILL44_32 VDD VSS sg13g2_FILL8
XSTDFILL44_40 VDD VSS sg13g2_FILL8
XSTDFILL44_48 VDD VSS sg13g2_FILL8
XSTDFILL44_56 VDD VSS sg13g2_FILL8
XSTDFILL44_64 VDD VSS sg13g2_FILL8
XSTDFILL44_72 VDD VSS sg13g2_FILL8
XSTDFILL44_80 VDD VSS sg13g2_FILL8
XSTDFILL44_88 VDD VSS sg13g2_FILL8
XSTDFILL44_96 VDD VSS sg13g2_FILL8
XSTDFILL44_104 VDD VSS sg13g2_FILL1
XSTDFILL44_1880 VDD VSS sg13g2_FILL8
XSTDFILL44_1888 VDD VSS sg13g2_FILL8
XSTDFILL44_1896 VDD VSS sg13g2_FILL8
XSTDFILL44_1904 VDD VSS sg13g2_FILL8
XSTDFILL44_1912 VDD VSS sg13g2_FILL8
XSTDFILL44_1920 VDD VSS sg13g2_FILL8
XSTDFILL44_1928 VDD VSS sg13g2_FILL8
XSTDFILL44_1936 VDD VSS sg13g2_FILL8
XSTDFILL44_1944 VDD VSS sg13g2_FILL8
XSTDFILL44_1952 VDD VSS sg13g2_FILL8
XSTDFILL44_1960 VDD VSS sg13g2_FILL8
XSTDFILL44_1968 VDD VSS sg13g2_FILL8
XSTDFILL44_1976 VDD VSS sg13g2_FILL8
XSTDFILL44_1984 VDD VSS sg13g2_FILL8
XSTDFILL44_1992 VDD VSS sg13g2_FILL8
XSTDFILL44_2000 VDD VSS sg13g2_FILL8
XSTDFILL44_2008 VDD VSS sg13g2_FILL8
XSTDFILL44_2016 VDD VSS sg13g2_FILL8
XSTDFILL44_2024 VDD VSS sg13g2_FILL8
XSTDFILL44_2032 VDD VSS sg13g2_FILL8
XSTDFILL44_2040 VDD VSS sg13g2_FILL8
XSTDFILL44_2048 VDD VSS sg13g2_FILL8
XSTDFILL44_2056 VDD VSS sg13g2_FILL8
XSTDFILL44_2064 VDD VSS sg13g2_FILL8
XSTDFILL44_2072 VDD VSS sg13g2_FILL8
XSTDFILL44_2080 VDD VSS sg13g2_FILL8
XSTDFILL44_2088 VDD VSS sg13g2_FILL8
XSTDFILL44_2096 VDD VSS sg13g2_FILL8
XSTDFILL44_2104 VDD VSS sg13g2_FILL8
XSTDFILL44_2112 VDD VSS sg13g2_FILL8
XSTDFILL44_2120 VDD VSS sg13g2_FILL8
XSTDFILL44_2128 VDD VSS sg13g2_FILL8
XSTDFILL44_2136 VDD VSS sg13g2_FILL8
XSTDFILL44_2144 VDD VSS sg13g2_FILL8
XSTDFILL44_2152 VDD VSS sg13g2_FILL8
XSTDFILL44_2160 VDD VSS sg13g2_FILL8
XSTDFILL44_2168 VDD VSS sg13g2_FILL4
XSTDFILL45_0 VDD VSS sg13g2_FILL8
XSTDFILL45_8 VDD VSS sg13g2_FILL8
XSTDFILL45_16 VDD VSS sg13g2_FILL8
XSTDFILL45_24 VDD VSS sg13g2_FILL8
XSTDFILL45_32 VDD VSS sg13g2_FILL8
XSTDFILL45_40 VDD VSS sg13g2_FILL8
XSTDFILL45_48 VDD VSS sg13g2_FILL8
XSTDFILL45_56 VDD VSS sg13g2_FILL8
XSTDFILL45_64 VDD VSS sg13g2_FILL8
XSTDFILL45_72 VDD VSS sg13g2_FILL8
XSTDFILL45_80 VDD VSS sg13g2_FILL8
XSTDFILL45_88 VDD VSS sg13g2_FILL8
XSTDFILL45_96 VDD VSS sg13g2_FILL8
XSTDFILL45_104 VDD VSS sg13g2_FILL1
XSTDFILL45_1880 VDD VSS sg13g2_FILL8
XSTDFILL45_1888 VDD VSS sg13g2_FILL8
XSTDFILL45_1896 VDD VSS sg13g2_FILL8
XSTDFILL45_1904 VDD VSS sg13g2_FILL8
XSTDFILL45_1912 VDD VSS sg13g2_FILL8
XSTDFILL45_1920 VDD VSS sg13g2_FILL8
XSTDFILL45_1928 VDD VSS sg13g2_FILL8
XSTDFILL45_1936 VDD VSS sg13g2_FILL8
XSTDFILL45_1944 VDD VSS sg13g2_FILL8
XSTDFILL45_1959 VDD VSS sg13g2_FILL8
XSTDFILL45_1967 VDD VSS sg13g2_FILL8
XSTDFILL45_1975 VDD VSS sg13g2_FILL8
XSTDFILL45_1983 VDD VSS sg13g2_FILL8
XSTDFILL45_1991 VDD VSS sg13g2_FILL4
XSTDFILL45_1995 VDD VSS sg13g2_FILL2
XSTDFILL45_1997 VDD VSS sg13g2_FILL1
XSTDFILL45_2005 VDD VSS sg13g2_FILL8
XSTDFILL45_2013 VDD VSS sg13g2_FILL8
XSTDFILL45_2021 VDD VSS sg13g2_FILL8
XSTDFILL45_2029 VDD VSS sg13g2_FILL8
XSTDFILL45_2037 VDD VSS sg13g2_FILL8
XSTDFILL45_2045 VDD VSS sg13g2_FILL8
XSTDFILL45_2053 VDD VSS sg13g2_FILL8
XSTDFILL45_2061 VDD VSS sg13g2_FILL8
XSTDFILL45_2069 VDD VSS sg13g2_FILL8
XSTDFILL45_2077 VDD VSS sg13g2_FILL8
XSTDFILL45_2085 VDD VSS sg13g2_FILL8
XSTDFILL45_2093 VDD VSS sg13g2_FILL8
XSTDFILL45_2101 VDD VSS sg13g2_FILL8
XSTDFILL45_2109 VDD VSS sg13g2_FILL8
XSTDFILL45_2117 VDD VSS sg13g2_FILL8
XSTDFILL45_2125 VDD VSS sg13g2_FILL8
XSTDFILL45_2133 VDD VSS sg13g2_FILL8
XSTDFILL45_2141 VDD VSS sg13g2_FILL8
XSTDFILL45_2149 VDD VSS sg13g2_FILL8
XSTDFILL45_2157 VDD VSS sg13g2_FILL8
XSTDFILL45_2165 VDD VSS sg13g2_FILL4
XSTDFILL45_2169 VDD VSS sg13g2_FILL2
XSTDFILL45_2171 VDD VSS sg13g2_FILL1
XSTDFILL46_0 VDD VSS sg13g2_FILL8
XSTDFILL46_8 VDD VSS sg13g2_FILL8
XSTDFILL46_16 VDD VSS sg13g2_FILL8
XSTDFILL46_24 VDD VSS sg13g2_FILL8
XSTDFILL46_32 VDD VSS sg13g2_FILL8
XSTDFILL46_40 VDD VSS sg13g2_FILL8
XSTDFILL46_48 VDD VSS sg13g2_FILL8
XSTDFILL46_56 VDD VSS sg13g2_FILL8
XSTDFILL46_64 VDD VSS sg13g2_FILL8
XSTDFILL46_72 VDD VSS sg13g2_FILL8
XSTDFILL46_80 VDD VSS sg13g2_FILL8
XSTDFILL46_88 VDD VSS sg13g2_FILL8
XSTDFILL46_96 VDD VSS sg13g2_FILL8
XSTDFILL46_104 VDD VSS sg13g2_FILL1
XSTDFILL46_1880 VDD VSS sg13g2_FILL8
XSTDFILL46_1888 VDD VSS sg13g2_FILL8
XSTDFILL46_1896 VDD VSS sg13g2_FILL8
XSTDFILL46_1904 VDD VSS sg13g2_FILL8
XSTDFILL46_1912 VDD VSS sg13g2_FILL8
XSTDFILL46_1920 VDD VSS sg13g2_FILL8
XSTDFILL46_1928 VDD VSS sg13g2_FILL8
XSTDFILL46_1936 VDD VSS sg13g2_FILL8
XSTDFILL46_1944 VDD VSS sg13g2_FILL1
XSTDFILL46_1960 VDD VSS sg13g2_FILL8
XSTDFILL46_1968 VDD VSS sg13g2_FILL8
XSTDFILL46_1976 VDD VSS sg13g2_FILL8
XSTDFILL46_1984 VDD VSS sg13g2_FILL4
XSTDFILL46_1988 VDD VSS sg13g2_FILL2
XSTDFILL46_1990 VDD VSS sg13g2_FILL1
XSTDFILL46_2006 VDD VSS sg13g2_FILL8
XSTDFILL46_2014 VDD VSS sg13g2_FILL8
XSTDFILL46_2022 VDD VSS sg13g2_FILL8
XSTDFILL46_2030 VDD VSS sg13g2_FILL8
XSTDFILL46_2038 VDD VSS sg13g2_FILL8
XSTDFILL46_2046 VDD VSS sg13g2_FILL8
XSTDFILL46_2054 VDD VSS sg13g2_FILL8
XSTDFILL46_2062 VDD VSS sg13g2_FILL8
XSTDFILL46_2070 VDD VSS sg13g2_FILL8
XSTDFILL46_2078 VDD VSS sg13g2_FILL8
XSTDFILL46_2086 VDD VSS sg13g2_FILL8
XSTDFILL46_2094 VDD VSS sg13g2_FILL8
XSTDFILL46_2102 VDD VSS sg13g2_FILL8
XSTDFILL46_2110 VDD VSS sg13g2_FILL8
XSTDFILL46_2118 VDD VSS sg13g2_FILL8
XSTDFILL46_2126 VDD VSS sg13g2_FILL8
XSTDFILL46_2134 VDD VSS sg13g2_FILL8
XSTDFILL46_2142 VDD VSS sg13g2_FILL8
XSTDFILL46_2150 VDD VSS sg13g2_FILL8
XSTDFILL46_2158 VDD VSS sg13g2_FILL8
XSTDFILL46_2166 VDD VSS sg13g2_FILL4
XSTDFILL46_2170 VDD VSS sg13g2_FILL2
XSTDFILL47_0 VDD VSS sg13g2_FILL8
XSTDFILL47_8 VDD VSS sg13g2_FILL8
XSTDFILL47_16 VDD VSS sg13g2_FILL8
XSTDFILL47_24 VDD VSS sg13g2_FILL8
XSTDFILL47_32 VDD VSS sg13g2_FILL8
XSTDFILL47_40 VDD VSS sg13g2_FILL8
XSTDFILL47_48 VDD VSS sg13g2_FILL8
XSTDFILL47_56 VDD VSS sg13g2_FILL8
XSTDFILL47_64 VDD VSS sg13g2_FILL8
XSTDFILL47_72 VDD VSS sg13g2_FILL8
XSTDFILL47_80 VDD VSS sg13g2_FILL8
XSTDFILL47_88 VDD VSS sg13g2_FILL8
XSTDFILL47_96 VDD VSS sg13g2_FILL8
XSTDFILL47_104 VDD VSS sg13g2_FILL1
XSTDFILL47_1880 VDD VSS sg13g2_FILL8
XSTDFILL47_1888 VDD VSS sg13g2_FILL8
XSTDFILL47_1896 VDD VSS sg13g2_FILL8
XSTDFILL47_1904 VDD VSS sg13g2_FILL8
XSTDFILL47_1912 VDD VSS sg13g2_FILL8
XSTDFILL47_1920 VDD VSS sg13g2_FILL8
XSTDFILL47_1928 VDD VSS sg13g2_FILL8
XSTDFILL47_1936 VDD VSS sg13g2_FILL8
XSTDFILL47_1944 VDD VSS sg13g2_FILL8
XSTDFILL47_1952 VDD VSS sg13g2_FILL8
XSTDFILL47_1960 VDD VSS sg13g2_FILL8
XSTDFILL47_1968 VDD VSS sg13g2_FILL8
XSTDFILL47_1976 VDD VSS sg13g2_FILL8
XSTDFILL47_1984 VDD VSS sg13g2_FILL8
XSTDFILL47_1992 VDD VSS sg13g2_FILL8
XSTDFILL47_2000 VDD VSS sg13g2_FILL8
XSTDFILL47_2008 VDD VSS sg13g2_FILL8
XSTDFILL47_2016 VDD VSS sg13g2_FILL8
XSTDFILL47_2024 VDD VSS sg13g2_FILL8
XSTDFILL47_2032 VDD VSS sg13g2_FILL8
XSTDFILL47_2040 VDD VSS sg13g2_FILL8
XSTDFILL47_2048 VDD VSS sg13g2_FILL8
XSTDFILL47_2056 VDD VSS sg13g2_FILL8
XSTDFILL47_2064 VDD VSS sg13g2_FILL8
XSTDFILL47_2072 VDD VSS sg13g2_FILL8
XSTDFILL47_2080 VDD VSS sg13g2_FILL8
XSTDFILL47_2088 VDD VSS sg13g2_FILL8
XSTDFILL47_2096 VDD VSS sg13g2_FILL8
XSTDFILL47_2104 VDD VSS sg13g2_FILL8
XSTDFILL47_2112 VDD VSS sg13g2_FILL8
XSTDFILL47_2120 VDD VSS sg13g2_FILL8
XSTDFILL47_2128 VDD VSS sg13g2_FILL8
XSTDFILL47_2136 VDD VSS sg13g2_FILL8
XSTDFILL47_2144 VDD VSS sg13g2_FILL8
XSTDFILL47_2152 VDD VSS sg13g2_FILL8
XSTDFILL47_2160 VDD VSS sg13g2_FILL8
XSTDFILL47_2168 VDD VSS sg13g2_FILL4
XSTDFILL48_0 VDD VSS sg13g2_FILL8
XSTDFILL48_8 VDD VSS sg13g2_FILL8
XSTDFILL48_16 VDD VSS sg13g2_FILL8
XSTDFILL48_24 VDD VSS sg13g2_FILL8
XSTDFILL48_32 VDD VSS sg13g2_FILL8
XSTDFILL48_40 VDD VSS sg13g2_FILL8
XSTDFILL48_48 VDD VSS sg13g2_FILL8
XSTDFILL48_56 VDD VSS sg13g2_FILL8
XSTDFILL48_64 VDD VSS sg13g2_FILL8
XSTDFILL48_72 VDD VSS sg13g2_FILL8
XSTDFILL48_80 VDD VSS sg13g2_FILL8
XSTDFILL48_88 VDD VSS sg13g2_FILL8
XSTDFILL48_96 VDD VSS sg13g2_FILL8
XSTDFILL48_104 VDD VSS sg13g2_FILL1
XSTDFILL48_1880 VDD VSS sg13g2_FILL8
XSTDFILL48_1888 VDD VSS sg13g2_FILL8
XSTDFILL48_1896 VDD VSS sg13g2_FILL8
XSTDFILL48_1904 VDD VSS sg13g2_FILL8
XSTDFILL48_1912 VDD VSS sg13g2_FILL8
XSTDFILL48_1920 VDD VSS sg13g2_FILL8
XSTDFILL48_1928 VDD VSS sg13g2_FILL8
XSTDFILL48_1936 VDD VSS sg13g2_FILL8
XSTDFILL48_1944 VDD VSS sg13g2_FILL8
XSTDFILL48_1952 VDD VSS sg13g2_FILL8
XSTDFILL48_1960 VDD VSS sg13g2_FILL8
XSTDFILL48_1968 VDD VSS sg13g2_FILL8
XSTDFILL48_1976 VDD VSS sg13g2_FILL8
XSTDFILL48_1984 VDD VSS sg13g2_FILL8
XSTDFILL48_1992 VDD VSS sg13g2_FILL8
XSTDFILL48_2000 VDD VSS sg13g2_FILL8
XSTDFILL48_2008 VDD VSS sg13g2_FILL8
XSTDFILL48_2016 VDD VSS sg13g2_FILL8
XSTDFILL48_2024 VDD VSS sg13g2_FILL8
XSTDFILL48_2032 VDD VSS sg13g2_FILL8
XSTDFILL48_2040 VDD VSS sg13g2_FILL8
XSTDFILL48_2048 VDD VSS sg13g2_FILL8
XSTDFILL48_2056 VDD VSS sg13g2_FILL8
XSTDFILL48_2064 VDD VSS sg13g2_FILL8
XSTDFILL48_2072 VDD VSS sg13g2_FILL8
XSTDFILL48_2080 VDD VSS sg13g2_FILL8
XSTDFILL48_2088 VDD VSS sg13g2_FILL8
XSTDFILL48_2096 VDD VSS sg13g2_FILL8
XSTDFILL48_2104 VDD VSS sg13g2_FILL8
XSTDFILL48_2112 VDD VSS sg13g2_FILL8
XSTDFILL48_2120 VDD VSS sg13g2_FILL8
XSTDFILL48_2128 VDD VSS sg13g2_FILL8
XSTDFILL48_2136 VDD VSS sg13g2_FILL8
XSTDFILL48_2144 VDD VSS sg13g2_FILL8
XSTDFILL48_2152 VDD VSS sg13g2_FILL8
XSTDFILL48_2160 VDD VSS sg13g2_FILL8
XSTDFILL48_2168 VDD VSS sg13g2_FILL4
XSTDFILL49_0 VDD VSS sg13g2_FILL8
XSTDFILL49_8 VDD VSS sg13g2_FILL8
XSTDFILL49_16 VDD VSS sg13g2_FILL8
XSTDFILL49_24 VDD VSS sg13g2_FILL8
XSTDFILL49_32 VDD VSS sg13g2_FILL8
XSTDFILL49_40 VDD VSS sg13g2_FILL8
XSTDFILL49_48 VDD VSS sg13g2_FILL8
XSTDFILL49_56 VDD VSS sg13g2_FILL8
XSTDFILL49_64 VDD VSS sg13g2_FILL8
XSTDFILL49_72 VDD VSS sg13g2_FILL8
XSTDFILL49_80 VDD VSS sg13g2_FILL8
XSTDFILL49_88 VDD VSS sg13g2_FILL8
XSTDFILL49_96 VDD VSS sg13g2_FILL8
XSTDFILL49_104 VDD VSS sg13g2_FILL1
XSTDFILL49_1880 VDD VSS sg13g2_FILL8
XSTDFILL49_1888 VDD VSS sg13g2_FILL8
XSTDFILL49_1896 VDD VSS sg13g2_FILL8
XSTDFILL49_1904 VDD VSS sg13g2_FILL8
XSTDFILL49_1912 VDD VSS sg13g2_FILL8
XSTDFILL49_1920 VDD VSS sg13g2_FILL8
XSTDFILL49_1928 VDD VSS sg13g2_FILL8
XSTDFILL49_1936 VDD VSS sg13g2_FILL8
XSTDFILL49_1944 VDD VSS sg13g2_FILL8
XSTDFILL49_1952 VDD VSS sg13g2_FILL8
XSTDFILL49_1960 VDD VSS sg13g2_FILL8
XSTDFILL49_1968 VDD VSS sg13g2_FILL8
XSTDFILL49_1976 VDD VSS sg13g2_FILL8
XSTDFILL49_1984 VDD VSS sg13g2_FILL8
XSTDFILL49_1992 VDD VSS sg13g2_FILL8
XSTDFILL49_2000 VDD VSS sg13g2_FILL8
XSTDFILL49_2008 VDD VSS sg13g2_FILL8
XSTDFILL49_2016 VDD VSS sg13g2_FILL8
XSTDFILL49_2024 VDD VSS sg13g2_FILL8
XSTDFILL49_2032 VDD VSS sg13g2_FILL8
XSTDFILL49_2040 VDD VSS sg13g2_FILL8
XSTDFILL49_2048 VDD VSS sg13g2_FILL8
XSTDFILL49_2056 VDD VSS sg13g2_FILL8
XSTDFILL49_2064 VDD VSS sg13g2_FILL8
XSTDFILL49_2072 VDD VSS sg13g2_FILL8
XSTDFILL49_2080 VDD VSS sg13g2_FILL8
XSTDFILL49_2088 VDD VSS sg13g2_FILL8
XSTDFILL49_2096 VDD VSS sg13g2_FILL8
XSTDFILL49_2104 VDD VSS sg13g2_FILL8
XSTDFILL49_2112 VDD VSS sg13g2_FILL8
XSTDFILL49_2120 VDD VSS sg13g2_FILL8
XSTDFILL49_2128 VDD VSS sg13g2_FILL8
XSTDFILL49_2136 VDD VSS sg13g2_FILL8
XSTDFILL49_2144 VDD VSS sg13g2_FILL8
XSTDFILL49_2152 VDD VSS sg13g2_FILL8
XSTDFILL49_2160 VDD VSS sg13g2_FILL8
XSTDFILL49_2168 VDD VSS sg13g2_FILL4
XSTDFILL50_0 VDD VSS sg13g2_FILL8
XSTDFILL50_8 VDD VSS sg13g2_FILL8
XSTDFILL50_16 VDD VSS sg13g2_FILL8
XSTDFILL50_24 VDD VSS sg13g2_FILL8
XSTDFILL50_32 VDD VSS sg13g2_FILL8
XSTDFILL50_40 VDD VSS sg13g2_FILL8
XSTDFILL50_48 VDD VSS sg13g2_FILL8
XSTDFILL50_56 VDD VSS sg13g2_FILL8
XSTDFILL50_64 VDD VSS sg13g2_FILL8
XSTDFILL50_72 VDD VSS sg13g2_FILL8
XSTDFILL50_80 VDD VSS sg13g2_FILL8
XSTDFILL50_88 VDD VSS sg13g2_FILL8
XSTDFILL50_96 VDD VSS sg13g2_FILL8
XSTDFILL50_104 VDD VSS sg13g2_FILL1
XSTDFILL50_1880 VDD VSS sg13g2_FILL8
XSTDFILL50_1888 VDD VSS sg13g2_FILL8
XSTDFILL50_1896 VDD VSS sg13g2_FILL8
XSTDFILL50_1904 VDD VSS sg13g2_FILL8
XSTDFILL50_1912 VDD VSS sg13g2_FILL8
XSTDFILL50_1920 VDD VSS sg13g2_FILL8
XSTDFILL50_1928 VDD VSS sg13g2_FILL8
XSTDFILL50_1936 VDD VSS sg13g2_FILL8
XSTDFILL50_1944 VDD VSS sg13g2_FILL8
XSTDFILL50_1952 VDD VSS sg13g2_FILL8
XSTDFILL50_1960 VDD VSS sg13g2_FILL8
XSTDFILL50_1968 VDD VSS sg13g2_FILL8
XSTDFILL50_1976 VDD VSS sg13g2_FILL8
XSTDFILL50_1984 VDD VSS sg13g2_FILL8
XSTDFILL50_1992 VDD VSS sg13g2_FILL8
XSTDFILL50_2000 VDD VSS sg13g2_FILL8
XSTDFILL50_2008 VDD VSS sg13g2_FILL8
XSTDFILL50_2016 VDD VSS sg13g2_FILL8
XSTDFILL50_2024 VDD VSS sg13g2_FILL8
XSTDFILL50_2032 VDD VSS sg13g2_FILL8
XSTDFILL50_2040 VDD VSS sg13g2_FILL8
XSTDFILL50_2048 VDD VSS sg13g2_FILL8
XSTDFILL50_2056 VDD VSS sg13g2_FILL8
XSTDFILL50_2064 VDD VSS sg13g2_FILL8
XSTDFILL50_2072 VDD VSS sg13g2_FILL8
XSTDFILL50_2080 VDD VSS sg13g2_FILL8
XSTDFILL50_2088 VDD VSS sg13g2_FILL8
XSTDFILL50_2096 VDD VSS sg13g2_FILL8
XSTDFILL50_2104 VDD VSS sg13g2_FILL8
XSTDFILL50_2112 VDD VSS sg13g2_FILL8
XSTDFILL50_2120 VDD VSS sg13g2_FILL8
XSTDFILL50_2128 VDD VSS sg13g2_FILL8
XSTDFILL50_2136 VDD VSS sg13g2_FILL8
XSTDFILL50_2144 VDD VSS sg13g2_FILL8
XSTDFILL50_2152 VDD VSS sg13g2_FILL8
XSTDFILL50_2160 VDD VSS sg13g2_FILL8
XSTDFILL50_2168 VDD VSS sg13g2_FILL4
XSTDFILL51_0 VDD VSS sg13g2_FILL8
XSTDFILL51_8 VDD VSS sg13g2_FILL8
XSTDFILL51_16 VDD VSS sg13g2_FILL8
XSTDFILL51_24 VDD VSS sg13g2_FILL8
XSTDFILL51_32 VDD VSS sg13g2_FILL8
XSTDFILL51_40 VDD VSS sg13g2_FILL8
XSTDFILL51_48 VDD VSS sg13g2_FILL8
XSTDFILL51_56 VDD VSS sg13g2_FILL8
XSTDFILL51_64 VDD VSS sg13g2_FILL8
XSTDFILL51_72 VDD VSS sg13g2_FILL8
XSTDFILL51_80 VDD VSS sg13g2_FILL8
XSTDFILL51_88 VDD VSS sg13g2_FILL8
XSTDFILL51_96 VDD VSS sg13g2_FILL8
XSTDFILL51_104 VDD VSS sg13g2_FILL1
XSTDFILL51_1880 VDD VSS sg13g2_FILL8
XSTDFILL51_1888 VDD VSS sg13g2_FILL8
XSTDFILL51_1896 VDD VSS sg13g2_FILL8
XSTDFILL51_1904 VDD VSS sg13g2_FILL8
XSTDFILL51_1912 VDD VSS sg13g2_FILL8
XSTDFILL51_1920 VDD VSS sg13g2_FILL8
XSTDFILL51_1928 VDD VSS sg13g2_FILL8
XSTDFILL51_1936 VDD VSS sg13g2_FILL8
XSTDFILL51_1944 VDD VSS sg13g2_FILL8
XSTDFILL51_1952 VDD VSS sg13g2_FILL8
XSTDFILL51_1960 VDD VSS sg13g2_FILL8
XSTDFILL51_1968 VDD VSS sg13g2_FILL8
XSTDFILL51_1976 VDD VSS sg13g2_FILL8
XSTDFILL51_1984 VDD VSS sg13g2_FILL8
XSTDFILL51_1992 VDD VSS sg13g2_FILL8
XSTDFILL51_2000 VDD VSS sg13g2_FILL8
XSTDFILL51_2008 VDD VSS sg13g2_FILL8
XSTDFILL51_2016 VDD VSS sg13g2_FILL8
XSTDFILL51_2024 VDD VSS sg13g2_FILL8
XSTDFILL51_2032 VDD VSS sg13g2_FILL8
XSTDFILL51_2040 VDD VSS sg13g2_FILL8
XSTDFILL51_2048 VDD VSS sg13g2_FILL8
XSTDFILL51_2056 VDD VSS sg13g2_FILL8
XSTDFILL51_2064 VDD VSS sg13g2_FILL8
XSTDFILL51_2072 VDD VSS sg13g2_FILL8
XSTDFILL51_2080 VDD VSS sg13g2_FILL8
XSTDFILL51_2088 VDD VSS sg13g2_FILL8
XSTDFILL51_2096 VDD VSS sg13g2_FILL8
XSTDFILL51_2104 VDD VSS sg13g2_FILL8
XSTDFILL51_2112 VDD VSS sg13g2_FILL8
XSTDFILL51_2120 VDD VSS sg13g2_FILL8
XSTDFILL51_2128 VDD VSS sg13g2_FILL8
XSTDFILL51_2136 VDD VSS sg13g2_FILL8
XSTDFILL51_2144 VDD VSS sg13g2_FILL8
XSTDFILL51_2152 VDD VSS sg13g2_FILL8
XSTDFILL51_2160 VDD VSS sg13g2_FILL8
XSTDFILL51_2168 VDD VSS sg13g2_FILL4
XSTDFILL52_0 VDD VSS sg13g2_FILL8
XSTDFILL52_8 VDD VSS sg13g2_FILL8
XSTDFILL52_16 VDD VSS sg13g2_FILL8
XSTDFILL52_24 VDD VSS sg13g2_FILL8
XSTDFILL52_32 VDD VSS sg13g2_FILL8
XSTDFILL52_40 VDD VSS sg13g2_FILL8
XSTDFILL52_48 VDD VSS sg13g2_FILL8
XSTDFILL52_56 VDD VSS sg13g2_FILL8
XSTDFILL52_64 VDD VSS sg13g2_FILL8
XSTDFILL52_72 VDD VSS sg13g2_FILL8
XSTDFILL52_80 VDD VSS sg13g2_FILL8
XSTDFILL52_88 VDD VSS sg13g2_FILL8
XSTDFILL52_96 VDD VSS sg13g2_FILL8
XSTDFILL52_104 VDD VSS sg13g2_FILL1
XSTDFILL52_1880 VDD VSS sg13g2_FILL8
XSTDFILL52_1888 VDD VSS sg13g2_FILL8
XSTDFILL52_1896 VDD VSS sg13g2_FILL8
XSTDFILL52_1904 VDD VSS sg13g2_FILL8
XSTDFILL52_1912 VDD VSS sg13g2_FILL8
XSTDFILL52_1920 VDD VSS sg13g2_FILL8
XSTDFILL52_1928 VDD VSS sg13g2_FILL8
XSTDFILL52_1936 VDD VSS sg13g2_FILL8
XSTDFILL52_1944 VDD VSS sg13g2_FILL8
XSTDFILL52_1952 VDD VSS sg13g2_FILL8
XSTDFILL52_1960 VDD VSS sg13g2_FILL8
XSTDFILL52_1968 VDD VSS sg13g2_FILL8
XSTDFILL52_1976 VDD VSS sg13g2_FILL8
XSTDFILL52_1984 VDD VSS sg13g2_FILL8
XSTDFILL52_1992 VDD VSS sg13g2_FILL8
XSTDFILL52_2000 VDD VSS sg13g2_FILL8
XSTDFILL52_2008 VDD VSS sg13g2_FILL8
XSTDFILL52_2016 VDD VSS sg13g2_FILL8
XSTDFILL52_2024 VDD VSS sg13g2_FILL8
XSTDFILL52_2032 VDD VSS sg13g2_FILL8
XSTDFILL52_2040 VDD VSS sg13g2_FILL8
XSTDFILL52_2048 VDD VSS sg13g2_FILL8
XSTDFILL52_2056 VDD VSS sg13g2_FILL8
XSTDFILL52_2064 VDD VSS sg13g2_FILL8
XSTDFILL52_2072 VDD VSS sg13g2_FILL8
XSTDFILL52_2080 VDD VSS sg13g2_FILL8
XSTDFILL52_2088 VDD VSS sg13g2_FILL8
XSTDFILL52_2096 VDD VSS sg13g2_FILL8
XSTDFILL52_2104 VDD VSS sg13g2_FILL8
XSTDFILL52_2112 VDD VSS sg13g2_FILL8
XSTDFILL52_2120 VDD VSS sg13g2_FILL8
XSTDFILL52_2128 VDD VSS sg13g2_FILL8
XSTDFILL52_2136 VDD VSS sg13g2_FILL8
XSTDFILL52_2144 VDD VSS sg13g2_FILL8
XSTDFILL52_2152 VDD VSS sg13g2_FILL8
XSTDFILL52_2160 VDD VSS sg13g2_FILL8
XSTDFILL52_2168 VDD VSS sg13g2_FILL4
XSTDFILL53_0 VDD VSS sg13g2_FILL8
XSTDFILL53_8 VDD VSS sg13g2_FILL8
XSTDFILL53_16 VDD VSS sg13g2_FILL8
XSTDFILL53_24 VDD VSS sg13g2_FILL8
XSTDFILL53_32 VDD VSS sg13g2_FILL8
XSTDFILL53_40 VDD VSS sg13g2_FILL8
XSTDFILL53_48 VDD VSS sg13g2_FILL8
XSTDFILL53_56 VDD VSS sg13g2_FILL8
XSTDFILL53_64 VDD VSS sg13g2_FILL8
XSTDFILL53_72 VDD VSS sg13g2_FILL8
XSTDFILL53_80 VDD VSS sg13g2_FILL8
XSTDFILL53_88 VDD VSS sg13g2_FILL8
XSTDFILL53_96 VDD VSS sg13g2_FILL8
XSTDFILL53_104 VDD VSS sg13g2_FILL1
XSTDFILL53_1880 VDD VSS sg13g2_FILL8
XSTDFILL53_1888 VDD VSS sg13g2_FILL8
XSTDFILL53_1896 VDD VSS sg13g2_FILL8
XSTDFILL53_1904 VDD VSS sg13g2_FILL8
XSTDFILL53_1912 VDD VSS sg13g2_FILL8
XSTDFILL53_1920 VDD VSS sg13g2_FILL8
XSTDFILL53_1928 VDD VSS sg13g2_FILL8
XSTDFILL53_1936 VDD VSS sg13g2_FILL8
XSTDFILL53_1944 VDD VSS sg13g2_FILL8
XSTDFILL53_1952 VDD VSS sg13g2_FILL8
XSTDFILL53_1960 VDD VSS sg13g2_FILL8
XSTDFILL53_1968 VDD VSS sg13g2_FILL8
XSTDFILL53_1976 VDD VSS sg13g2_FILL8
XSTDFILL53_1984 VDD VSS sg13g2_FILL8
XSTDFILL53_1992 VDD VSS sg13g2_FILL8
XSTDFILL53_2000 VDD VSS sg13g2_FILL8
XSTDFILL53_2008 VDD VSS sg13g2_FILL8
XSTDFILL53_2016 VDD VSS sg13g2_FILL8
XSTDFILL53_2024 VDD VSS sg13g2_FILL8
XSTDFILL53_2032 VDD VSS sg13g2_FILL8
XSTDFILL53_2040 VDD VSS sg13g2_FILL8
XSTDFILL53_2048 VDD VSS sg13g2_FILL8
XSTDFILL53_2056 VDD VSS sg13g2_FILL8
XSTDFILL53_2064 VDD VSS sg13g2_FILL8
XSTDFILL53_2072 VDD VSS sg13g2_FILL8
XSTDFILL53_2080 VDD VSS sg13g2_FILL8
XSTDFILL53_2088 VDD VSS sg13g2_FILL8
XSTDFILL53_2096 VDD VSS sg13g2_FILL8
XSTDFILL53_2104 VDD VSS sg13g2_FILL8
XSTDFILL53_2112 VDD VSS sg13g2_FILL8
XSTDFILL53_2120 VDD VSS sg13g2_FILL8
XSTDFILL53_2128 VDD VSS sg13g2_FILL8
XSTDFILL53_2136 VDD VSS sg13g2_FILL8
XSTDFILL53_2144 VDD VSS sg13g2_FILL8
XSTDFILL53_2152 VDD VSS sg13g2_FILL8
XSTDFILL53_2160 VDD VSS sg13g2_FILL8
XSTDFILL53_2168 VDD VSS sg13g2_FILL4
XSTDFILL54_0 VDD VSS sg13g2_FILL8
XSTDFILL54_8 VDD VSS sg13g2_FILL8
XSTDFILL54_16 VDD VSS sg13g2_FILL8
XSTDFILL54_24 VDD VSS sg13g2_FILL8
XSTDFILL54_32 VDD VSS sg13g2_FILL8
XSTDFILL54_40 VDD VSS sg13g2_FILL8
XSTDFILL54_48 VDD VSS sg13g2_FILL8
XSTDFILL54_56 VDD VSS sg13g2_FILL8
XSTDFILL54_64 VDD VSS sg13g2_FILL8
XSTDFILL54_72 VDD VSS sg13g2_FILL8
XSTDFILL54_80 VDD VSS sg13g2_FILL8
XSTDFILL54_88 VDD VSS sg13g2_FILL8
XSTDFILL54_96 VDD VSS sg13g2_FILL8
XSTDFILL54_104 VDD VSS sg13g2_FILL1
XSTDFILL54_1880 VDD VSS sg13g2_FILL8
XSTDFILL54_1888 VDD VSS sg13g2_FILL8
XSTDFILL54_1896 VDD VSS sg13g2_FILL8
XSTDFILL54_1904 VDD VSS sg13g2_FILL8
XSTDFILL54_1912 VDD VSS sg13g2_FILL8
XSTDFILL54_1920 VDD VSS sg13g2_FILL8
XSTDFILL54_1928 VDD VSS sg13g2_FILL8
XSTDFILL54_1936 VDD VSS sg13g2_FILL8
XSTDFILL54_1944 VDD VSS sg13g2_FILL8
XSTDFILL54_1952 VDD VSS sg13g2_FILL8
XSTDFILL54_1960 VDD VSS sg13g2_FILL8
XSTDFILL54_1968 VDD VSS sg13g2_FILL8
XSTDFILL54_1976 VDD VSS sg13g2_FILL8
XSTDFILL54_1984 VDD VSS sg13g2_FILL8
XSTDFILL54_1992 VDD VSS sg13g2_FILL8
XSTDFILL54_2000 VDD VSS sg13g2_FILL8
XSTDFILL54_2008 VDD VSS sg13g2_FILL8
XSTDFILL54_2016 VDD VSS sg13g2_FILL8
XSTDFILL54_2024 VDD VSS sg13g2_FILL8
XSTDFILL54_2032 VDD VSS sg13g2_FILL8
XSTDFILL54_2040 VDD VSS sg13g2_FILL8
XSTDFILL54_2048 VDD VSS sg13g2_FILL8
XSTDFILL54_2056 VDD VSS sg13g2_FILL8
XSTDFILL54_2064 VDD VSS sg13g2_FILL8
XSTDFILL54_2072 VDD VSS sg13g2_FILL8
XSTDFILL54_2080 VDD VSS sg13g2_FILL8
XSTDFILL54_2088 VDD VSS sg13g2_FILL8
XSTDFILL54_2096 VDD VSS sg13g2_FILL8
XSTDFILL54_2104 VDD VSS sg13g2_FILL8
XSTDFILL54_2112 VDD VSS sg13g2_FILL8
XSTDFILL54_2120 VDD VSS sg13g2_FILL8
XSTDFILL54_2128 VDD VSS sg13g2_FILL8
XSTDFILL54_2136 VDD VSS sg13g2_FILL8
XSTDFILL54_2144 VDD VSS sg13g2_FILL8
XSTDFILL54_2152 VDD VSS sg13g2_FILL8
XSTDFILL54_2160 VDD VSS sg13g2_FILL8
XSTDFILL54_2168 VDD VSS sg13g2_FILL4
XSTDFILL55_0 VDD VSS sg13g2_FILL8
XSTDFILL55_8 VDD VSS sg13g2_FILL8
XSTDFILL55_16 VDD VSS sg13g2_FILL8
XSTDFILL55_24 VDD VSS sg13g2_FILL8
XSTDFILL55_32 VDD VSS sg13g2_FILL8
XSTDFILL55_40 VDD VSS sg13g2_FILL8
XSTDFILL55_48 VDD VSS sg13g2_FILL8
XSTDFILL55_56 VDD VSS sg13g2_FILL8
XSTDFILL55_64 VDD VSS sg13g2_FILL8
XSTDFILL55_72 VDD VSS sg13g2_FILL8
XSTDFILL55_80 VDD VSS sg13g2_FILL8
XSTDFILL55_88 VDD VSS sg13g2_FILL8
XSTDFILL55_96 VDD VSS sg13g2_FILL8
XSTDFILL55_104 VDD VSS sg13g2_FILL1
XSTDFILL55_1880 VDD VSS sg13g2_FILL8
XSTDFILL55_1888 VDD VSS sg13g2_FILL8
XSTDFILL55_1896 VDD VSS sg13g2_FILL8
XSTDFILL55_1904 VDD VSS sg13g2_FILL8
XSTDFILL55_1912 VDD VSS sg13g2_FILL8
XSTDFILL55_1920 VDD VSS sg13g2_FILL8
XSTDFILL55_1928 VDD VSS sg13g2_FILL8
XSTDFILL55_1936 VDD VSS sg13g2_FILL8
XSTDFILL55_1944 VDD VSS sg13g2_FILL8
XSTDFILL55_1952 VDD VSS sg13g2_FILL8
XSTDFILL55_1960 VDD VSS sg13g2_FILL8
XSTDFILL55_1968 VDD VSS sg13g2_FILL8
XSTDFILL55_1976 VDD VSS sg13g2_FILL8
XSTDFILL55_1984 VDD VSS sg13g2_FILL8
XSTDFILL55_1992 VDD VSS sg13g2_FILL8
XSTDFILL55_2000 VDD VSS sg13g2_FILL8
XSTDFILL55_2008 VDD VSS sg13g2_FILL8
XSTDFILL55_2016 VDD VSS sg13g2_FILL8
XSTDFILL55_2024 VDD VSS sg13g2_FILL8
XSTDFILL55_2032 VDD VSS sg13g2_FILL8
XSTDFILL55_2040 VDD VSS sg13g2_FILL8
XSTDFILL55_2048 VDD VSS sg13g2_FILL8
XSTDFILL55_2056 VDD VSS sg13g2_FILL8
XSTDFILL55_2064 VDD VSS sg13g2_FILL8
XSTDFILL55_2072 VDD VSS sg13g2_FILL8
XSTDFILL55_2080 VDD VSS sg13g2_FILL8
XSTDFILL55_2088 VDD VSS sg13g2_FILL8
XSTDFILL55_2096 VDD VSS sg13g2_FILL8
XSTDFILL55_2104 VDD VSS sg13g2_FILL8
XSTDFILL55_2112 VDD VSS sg13g2_FILL8
XSTDFILL55_2120 VDD VSS sg13g2_FILL8
XSTDFILL55_2128 VDD VSS sg13g2_FILL8
XSTDFILL55_2136 VDD VSS sg13g2_FILL8
XSTDFILL55_2144 VDD VSS sg13g2_FILL8
XSTDFILL55_2152 VDD VSS sg13g2_FILL8
XSTDFILL55_2160 VDD VSS sg13g2_FILL8
XSTDFILL55_2168 VDD VSS sg13g2_FILL4
XSTDFILL56_0 VDD VSS sg13g2_FILL8
XSTDFILL56_8 VDD VSS sg13g2_FILL8
XSTDFILL56_16 VDD VSS sg13g2_FILL8
XSTDFILL56_24 VDD VSS sg13g2_FILL8
XSTDFILL56_32 VDD VSS sg13g2_FILL8
XSTDFILL56_40 VDD VSS sg13g2_FILL8
XSTDFILL56_48 VDD VSS sg13g2_FILL8
XSTDFILL56_56 VDD VSS sg13g2_FILL8
XSTDFILL56_64 VDD VSS sg13g2_FILL8
XSTDFILL56_72 VDD VSS sg13g2_FILL8
XSTDFILL56_80 VDD VSS sg13g2_FILL8
XSTDFILL56_88 VDD VSS sg13g2_FILL8
XSTDFILL56_96 VDD VSS sg13g2_FILL8
XSTDFILL56_104 VDD VSS sg13g2_FILL1
XSTDFILL56_1880 VDD VSS sg13g2_FILL8
XSTDFILL56_1888 VDD VSS sg13g2_FILL8
XSTDFILL56_1896 VDD VSS sg13g2_FILL8
XSTDFILL56_1904 VDD VSS sg13g2_FILL8
XSTDFILL56_1912 VDD VSS sg13g2_FILL8
XSTDFILL56_1920 VDD VSS sg13g2_FILL8
XSTDFILL56_1928 VDD VSS sg13g2_FILL8
XSTDFILL56_1936 VDD VSS sg13g2_FILL8
XSTDFILL56_1944 VDD VSS sg13g2_FILL8
XSTDFILL56_1952 VDD VSS sg13g2_FILL8
XSTDFILL56_1960 VDD VSS sg13g2_FILL8
XSTDFILL56_1968 VDD VSS sg13g2_FILL8
XSTDFILL56_1976 VDD VSS sg13g2_FILL8
XSTDFILL56_1984 VDD VSS sg13g2_FILL8
XSTDFILL56_1992 VDD VSS sg13g2_FILL8
XSTDFILL56_2000 VDD VSS sg13g2_FILL8
XSTDFILL56_2008 VDD VSS sg13g2_FILL8
XSTDFILL56_2016 VDD VSS sg13g2_FILL8
XSTDFILL56_2024 VDD VSS sg13g2_FILL8
XSTDFILL56_2032 VDD VSS sg13g2_FILL8
XSTDFILL56_2040 VDD VSS sg13g2_FILL8
XSTDFILL56_2048 VDD VSS sg13g2_FILL8
XSTDFILL56_2056 VDD VSS sg13g2_FILL8
XSTDFILL56_2064 VDD VSS sg13g2_FILL8
XSTDFILL56_2072 VDD VSS sg13g2_FILL8
XSTDFILL56_2080 VDD VSS sg13g2_FILL8
XSTDFILL56_2088 VDD VSS sg13g2_FILL8
XSTDFILL56_2096 VDD VSS sg13g2_FILL8
XSTDFILL56_2104 VDD VSS sg13g2_FILL8
XSTDFILL56_2112 VDD VSS sg13g2_FILL8
XSTDFILL56_2120 VDD VSS sg13g2_FILL8
XSTDFILL56_2128 VDD VSS sg13g2_FILL8
XSTDFILL56_2136 VDD VSS sg13g2_FILL8
XSTDFILL56_2144 VDD VSS sg13g2_FILL8
XSTDFILL56_2152 VDD VSS sg13g2_FILL8
XSTDFILL56_2160 VDD VSS sg13g2_FILL8
XSTDFILL56_2168 VDD VSS sg13g2_FILL4
XSTDFILL57_0 VDD VSS sg13g2_FILL8
XSTDFILL57_8 VDD VSS sg13g2_FILL8
XSTDFILL57_16 VDD VSS sg13g2_FILL8
XSTDFILL57_24 VDD VSS sg13g2_FILL8
XSTDFILL57_32 VDD VSS sg13g2_FILL8
XSTDFILL57_40 VDD VSS sg13g2_FILL8
XSTDFILL57_48 VDD VSS sg13g2_FILL8
XSTDFILL57_56 VDD VSS sg13g2_FILL8
XSTDFILL57_64 VDD VSS sg13g2_FILL8
XSTDFILL57_72 VDD VSS sg13g2_FILL8
XSTDFILL57_80 VDD VSS sg13g2_FILL8
XSTDFILL57_88 VDD VSS sg13g2_FILL8
XSTDFILL57_96 VDD VSS sg13g2_FILL8
XSTDFILL57_104 VDD VSS sg13g2_FILL1
XSTDFILL57_1880 VDD VSS sg13g2_FILL8
XSTDFILL57_1888 VDD VSS sg13g2_FILL8
XSTDFILL57_1896 VDD VSS sg13g2_FILL8
XSTDFILL57_1904 VDD VSS sg13g2_FILL8
XSTDFILL57_1912 VDD VSS sg13g2_FILL8
XSTDFILL57_1920 VDD VSS sg13g2_FILL8
XSTDFILL57_1928 VDD VSS sg13g2_FILL8
XSTDFILL57_1936 VDD VSS sg13g2_FILL8
XSTDFILL57_1944 VDD VSS sg13g2_FILL8
XSTDFILL57_1952 VDD VSS sg13g2_FILL8
XSTDFILL57_1960 VDD VSS sg13g2_FILL8
XSTDFILL57_1968 VDD VSS sg13g2_FILL8
XSTDFILL57_1976 VDD VSS sg13g2_FILL8
XSTDFILL57_1984 VDD VSS sg13g2_FILL8
XSTDFILL57_1992 VDD VSS sg13g2_FILL8
XSTDFILL57_2000 VDD VSS sg13g2_FILL8
XSTDFILL57_2008 VDD VSS sg13g2_FILL8
XSTDFILL57_2016 VDD VSS sg13g2_FILL8
XSTDFILL57_2024 VDD VSS sg13g2_FILL8
XSTDFILL57_2032 VDD VSS sg13g2_FILL8
XSTDFILL57_2040 VDD VSS sg13g2_FILL8
XSTDFILL57_2048 VDD VSS sg13g2_FILL8
XSTDFILL57_2056 VDD VSS sg13g2_FILL8
XSTDFILL57_2064 VDD VSS sg13g2_FILL8
XSTDFILL57_2072 VDD VSS sg13g2_FILL8
XSTDFILL57_2080 VDD VSS sg13g2_FILL8
XSTDFILL57_2088 VDD VSS sg13g2_FILL8
XSTDFILL57_2096 VDD VSS sg13g2_FILL8
XSTDFILL57_2104 VDD VSS sg13g2_FILL8
XSTDFILL57_2112 VDD VSS sg13g2_FILL8
XSTDFILL57_2120 VDD VSS sg13g2_FILL8
XSTDFILL57_2128 VDD VSS sg13g2_FILL8
XSTDFILL57_2136 VDD VSS sg13g2_FILL8
XSTDFILL57_2144 VDD VSS sg13g2_FILL8
XSTDFILL57_2152 VDD VSS sg13g2_FILL8
XSTDFILL57_2160 VDD VSS sg13g2_FILL8
XSTDFILL57_2168 VDD VSS sg13g2_FILL4
XSTDFILL58_0 VDD VSS sg13g2_FILL8
XSTDFILL58_8 VDD VSS sg13g2_FILL8
XSTDFILL58_16 VDD VSS sg13g2_FILL8
XSTDFILL58_24 VDD VSS sg13g2_FILL8
XSTDFILL58_32 VDD VSS sg13g2_FILL8
XSTDFILL58_40 VDD VSS sg13g2_FILL8
XSTDFILL58_48 VDD VSS sg13g2_FILL8
XSTDFILL58_56 VDD VSS sg13g2_FILL8
XSTDFILL58_64 VDD VSS sg13g2_FILL8
XSTDFILL58_72 VDD VSS sg13g2_FILL8
XSTDFILL58_80 VDD VSS sg13g2_FILL8
XSTDFILL58_88 VDD VSS sg13g2_FILL8
XSTDFILL58_96 VDD VSS sg13g2_FILL8
XSTDFILL58_104 VDD VSS sg13g2_FILL1
XSTDFILL58_1880 VDD VSS sg13g2_FILL8
XSTDFILL58_1888 VDD VSS sg13g2_FILL8
XSTDFILL58_1896 VDD VSS sg13g2_FILL8
XSTDFILL58_1904 VDD VSS sg13g2_FILL8
XSTDFILL58_1912 VDD VSS sg13g2_FILL8
XSTDFILL58_1920 VDD VSS sg13g2_FILL8
XSTDFILL58_1928 VDD VSS sg13g2_FILL8
XSTDFILL58_1936 VDD VSS sg13g2_FILL8
XSTDFILL58_1944 VDD VSS sg13g2_FILL8
XSTDFILL58_1952 VDD VSS sg13g2_FILL8
XSTDFILL58_1960 VDD VSS sg13g2_FILL8
XSTDFILL58_1968 VDD VSS sg13g2_FILL8
XSTDFILL58_1976 VDD VSS sg13g2_FILL8
XSTDFILL58_1984 VDD VSS sg13g2_FILL8
XSTDFILL58_1992 VDD VSS sg13g2_FILL8
XSTDFILL58_2000 VDD VSS sg13g2_FILL8
XSTDFILL58_2008 VDD VSS sg13g2_FILL8
XSTDFILL58_2016 VDD VSS sg13g2_FILL8
XSTDFILL58_2024 VDD VSS sg13g2_FILL8
XSTDFILL58_2032 VDD VSS sg13g2_FILL8
XSTDFILL58_2040 VDD VSS sg13g2_FILL8
XSTDFILL58_2048 VDD VSS sg13g2_FILL8
XSTDFILL58_2056 VDD VSS sg13g2_FILL8
XSTDFILL58_2064 VDD VSS sg13g2_FILL8
XSTDFILL58_2072 VDD VSS sg13g2_FILL8
XSTDFILL58_2080 VDD VSS sg13g2_FILL8
XSTDFILL58_2088 VDD VSS sg13g2_FILL8
XSTDFILL58_2096 VDD VSS sg13g2_FILL8
XSTDFILL58_2104 VDD VSS sg13g2_FILL8
XSTDFILL58_2112 VDD VSS sg13g2_FILL8
XSTDFILL58_2120 VDD VSS sg13g2_FILL8
XSTDFILL58_2128 VDD VSS sg13g2_FILL8
XSTDFILL58_2136 VDD VSS sg13g2_FILL8
XSTDFILL58_2144 VDD VSS sg13g2_FILL8
XSTDFILL58_2152 VDD VSS sg13g2_FILL8
XSTDFILL58_2160 VDD VSS sg13g2_FILL8
XSTDFILL58_2168 VDD VSS sg13g2_FILL4
XSTDFILL59_0 VDD VSS sg13g2_FILL8
XSTDFILL59_8 VDD VSS sg13g2_FILL8
XSTDFILL59_16 VDD VSS sg13g2_FILL8
XSTDFILL59_24 VDD VSS sg13g2_FILL8
XSTDFILL59_32 VDD VSS sg13g2_FILL8
XSTDFILL59_40 VDD VSS sg13g2_FILL8
XSTDFILL59_48 VDD VSS sg13g2_FILL8
XSTDFILL59_56 VDD VSS sg13g2_FILL8
XSTDFILL59_64 VDD VSS sg13g2_FILL8
XSTDFILL59_72 VDD VSS sg13g2_FILL8
XSTDFILL59_80 VDD VSS sg13g2_FILL8
XSTDFILL59_88 VDD VSS sg13g2_FILL8
XSTDFILL59_96 VDD VSS sg13g2_FILL8
XSTDFILL59_104 VDD VSS sg13g2_FILL1
XSTDFILL59_1880 VDD VSS sg13g2_FILL8
XSTDFILL59_1888 VDD VSS sg13g2_FILL8
XSTDFILL59_1896 VDD VSS sg13g2_FILL8
XSTDFILL59_1904 VDD VSS sg13g2_FILL8
XSTDFILL59_1912 VDD VSS sg13g2_FILL8
XSTDFILL59_1920 VDD VSS sg13g2_FILL8
XSTDFILL59_1928 VDD VSS sg13g2_FILL8
XSTDFILL59_1936 VDD VSS sg13g2_FILL8
XSTDFILL59_1944 VDD VSS sg13g2_FILL8
XSTDFILL59_1952 VDD VSS sg13g2_FILL8
XSTDFILL59_1960 VDD VSS sg13g2_FILL8
XSTDFILL59_1968 VDD VSS sg13g2_FILL8
XSTDFILL59_1976 VDD VSS sg13g2_FILL8
XSTDFILL59_1984 VDD VSS sg13g2_FILL8
XSTDFILL59_1992 VDD VSS sg13g2_FILL8
XSTDFILL59_2000 VDD VSS sg13g2_FILL8
XSTDFILL59_2008 VDD VSS sg13g2_FILL8
XSTDFILL59_2016 VDD VSS sg13g2_FILL8
XSTDFILL59_2024 VDD VSS sg13g2_FILL8
XSTDFILL59_2032 VDD VSS sg13g2_FILL8
XSTDFILL59_2040 VDD VSS sg13g2_FILL8
XSTDFILL59_2048 VDD VSS sg13g2_FILL8
XSTDFILL59_2056 VDD VSS sg13g2_FILL8
XSTDFILL59_2064 VDD VSS sg13g2_FILL8
XSTDFILL59_2072 VDD VSS sg13g2_FILL8
XSTDFILL59_2080 VDD VSS sg13g2_FILL8
XSTDFILL59_2088 VDD VSS sg13g2_FILL8
XSTDFILL59_2096 VDD VSS sg13g2_FILL8
XSTDFILL59_2104 VDD VSS sg13g2_FILL8
XSTDFILL59_2112 VDD VSS sg13g2_FILL8
XSTDFILL59_2120 VDD VSS sg13g2_FILL8
XSTDFILL59_2128 VDD VSS sg13g2_FILL8
XSTDFILL59_2136 VDD VSS sg13g2_FILL8
XSTDFILL59_2144 VDD VSS sg13g2_FILL8
XSTDFILL59_2152 VDD VSS sg13g2_FILL8
XSTDFILL59_2160 VDD VSS sg13g2_FILL8
XSTDFILL59_2168 VDD VSS sg13g2_FILL4
XSTDFILL60_0 VDD VSS sg13g2_FILL8
XSTDFILL60_8 VDD VSS sg13g2_FILL8
XSTDFILL60_16 VDD VSS sg13g2_FILL8
XSTDFILL60_24 VDD VSS sg13g2_FILL8
XSTDFILL60_32 VDD VSS sg13g2_FILL8
XSTDFILL60_40 VDD VSS sg13g2_FILL8
XSTDFILL60_48 VDD VSS sg13g2_FILL8
XSTDFILL60_56 VDD VSS sg13g2_FILL8
XSTDFILL60_64 VDD VSS sg13g2_FILL8
XSTDFILL60_72 VDD VSS sg13g2_FILL8
XSTDFILL60_80 VDD VSS sg13g2_FILL8
XSTDFILL60_88 VDD VSS sg13g2_FILL8
XSTDFILL60_96 VDD VSS sg13g2_FILL8
XSTDFILL60_104 VDD VSS sg13g2_FILL1
XSTDFILL60_1880 VDD VSS sg13g2_FILL8
XSTDFILL60_1888 VDD VSS sg13g2_FILL8
XSTDFILL60_1896 VDD VSS sg13g2_FILL8
XSTDFILL60_1904 VDD VSS sg13g2_FILL8
XSTDFILL60_1912 VDD VSS sg13g2_FILL8
XSTDFILL60_1920 VDD VSS sg13g2_FILL8
XSTDFILL60_1928 VDD VSS sg13g2_FILL8
XSTDFILL60_1936 VDD VSS sg13g2_FILL8
XSTDFILL60_1944 VDD VSS sg13g2_FILL8
XSTDFILL60_1952 VDD VSS sg13g2_FILL8
XSTDFILL60_1960 VDD VSS sg13g2_FILL8
XSTDFILL60_1968 VDD VSS sg13g2_FILL8
XSTDFILL60_1976 VDD VSS sg13g2_FILL8
XSTDFILL60_1984 VDD VSS sg13g2_FILL8
XSTDFILL60_1992 VDD VSS sg13g2_FILL8
XSTDFILL60_2000 VDD VSS sg13g2_FILL8
XSTDFILL60_2008 VDD VSS sg13g2_FILL8
XSTDFILL60_2016 VDD VSS sg13g2_FILL8
XSTDFILL60_2024 VDD VSS sg13g2_FILL8
XSTDFILL60_2032 VDD VSS sg13g2_FILL8
XSTDFILL60_2040 VDD VSS sg13g2_FILL8
XSTDFILL60_2048 VDD VSS sg13g2_FILL8
XSTDFILL60_2056 VDD VSS sg13g2_FILL8
XSTDFILL60_2064 VDD VSS sg13g2_FILL8
XSTDFILL60_2072 VDD VSS sg13g2_FILL8
XSTDFILL60_2080 VDD VSS sg13g2_FILL8
XSTDFILL60_2088 VDD VSS sg13g2_FILL8
XSTDFILL60_2096 VDD VSS sg13g2_FILL8
XSTDFILL60_2104 VDD VSS sg13g2_FILL8
XSTDFILL60_2112 VDD VSS sg13g2_FILL8
XSTDFILL60_2120 VDD VSS sg13g2_FILL8
XSTDFILL60_2128 VDD VSS sg13g2_FILL8
XSTDFILL60_2136 VDD VSS sg13g2_FILL8
XSTDFILL60_2144 VDD VSS sg13g2_FILL8
XSTDFILL60_2152 VDD VSS sg13g2_FILL8
XSTDFILL60_2160 VDD VSS sg13g2_FILL8
XSTDFILL60_2168 VDD VSS sg13g2_FILL4
XSTDFILL61_0 VDD VSS sg13g2_FILL8
XSTDFILL61_8 VDD VSS sg13g2_FILL8
XSTDFILL61_16 VDD VSS sg13g2_FILL8
XSTDFILL61_24 VDD VSS sg13g2_FILL8
XSTDFILL61_32 VDD VSS sg13g2_FILL8
XSTDFILL61_40 VDD VSS sg13g2_FILL8
XSTDFILL61_48 VDD VSS sg13g2_FILL8
XSTDFILL61_56 VDD VSS sg13g2_FILL8
XSTDFILL61_64 VDD VSS sg13g2_FILL8
XSTDFILL61_72 VDD VSS sg13g2_FILL8
XSTDFILL61_80 VDD VSS sg13g2_FILL8
XSTDFILL61_88 VDD VSS sg13g2_FILL8
XSTDFILL61_96 VDD VSS sg13g2_FILL8
XSTDFILL61_104 VDD VSS sg13g2_FILL1
XSTDFILL61_1880 VDD VSS sg13g2_FILL8
XSTDFILL61_1888 VDD VSS sg13g2_FILL8
XSTDFILL61_1896 VDD VSS sg13g2_FILL8
XSTDFILL61_1904 VDD VSS sg13g2_FILL8
XSTDFILL61_1912 VDD VSS sg13g2_FILL8
XSTDFILL61_1920 VDD VSS sg13g2_FILL8
XSTDFILL61_1928 VDD VSS sg13g2_FILL8
XSTDFILL61_1936 VDD VSS sg13g2_FILL8
XSTDFILL61_1944 VDD VSS sg13g2_FILL8
XSTDFILL61_1952 VDD VSS sg13g2_FILL8
XSTDFILL61_1960 VDD VSS sg13g2_FILL8
XSTDFILL61_1968 VDD VSS sg13g2_FILL8
XSTDFILL61_1976 VDD VSS sg13g2_FILL8
XSTDFILL61_1984 VDD VSS sg13g2_FILL8
XSTDFILL61_1992 VDD VSS sg13g2_FILL8
XSTDFILL61_2000 VDD VSS sg13g2_FILL8
XSTDFILL61_2008 VDD VSS sg13g2_FILL8
XSTDFILL61_2016 VDD VSS sg13g2_FILL8
XSTDFILL61_2024 VDD VSS sg13g2_FILL8
XSTDFILL61_2032 VDD VSS sg13g2_FILL8
XSTDFILL61_2040 VDD VSS sg13g2_FILL8
XSTDFILL61_2048 VDD VSS sg13g2_FILL8
XSTDFILL61_2056 VDD VSS sg13g2_FILL8
XSTDFILL61_2064 VDD VSS sg13g2_FILL8
XSTDFILL61_2072 VDD VSS sg13g2_FILL8
XSTDFILL61_2080 VDD VSS sg13g2_FILL8
XSTDFILL61_2088 VDD VSS sg13g2_FILL8
XSTDFILL61_2096 VDD VSS sg13g2_FILL8
XSTDFILL61_2104 VDD VSS sg13g2_FILL8
XSTDFILL61_2112 VDD VSS sg13g2_FILL8
XSTDFILL61_2120 VDD VSS sg13g2_FILL8
XSTDFILL61_2128 VDD VSS sg13g2_FILL8
XSTDFILL61_2136 VDD VSS sg13g2_FILL8
XSTDFILL61_2144 VDD VSS sg13g2_FILL8
XSTDFILL61_2152 VDD VSS sg13g2_FILL8
XSTDFILL61_2160 VDD VSS sg13g2_FILL8
XSTDFILL61_2168 VDD VSS sg13g2_FILL4
XSTDFILL62_0 VDD VSS sg13g2_FILL8
XSTDFILL62_8 VDD VSS sg13g2_FILL8
XSTDFILL62_16 VDD VSS sg13g2_FILL8
XSTDFILL62_24 VDD VSS sg13g2_FILL8
XSTDFILL62_32 VDD VSS sg13g2_FILL8
XSTDFILL62_40 VDD VSS sg13g2_FILL8
XSTDFILL62_48 VDD VSS sg13g2_FILL8
XSTDFILL62_56 VDD VSS sg13g2_FILL8
XSTDFILL62_64 VDD VSS sg13g2_FILL8
XSTDFILL62_72 VDD VSS sg13g2_FILL8
XSTDFILL62_80 VDD VSS sg13g2_FILL8
XSTDFILL62_88 VDD VSS sg13g2_FILL8
XSTDFILL62_96 VDD VSS sg13g2_FILL8
XSTDFILL62_104 VDD VSS sg13g2_FILL1
XSTDFILL62_1880 VDD VSS sg13g2_FILL8
XSTDFILL62_1888 VDD VSS sg13g2_FILL8
XSTDFILL62_1896 VDD VSS sg13g2_FILL8
XSTDFILL62_1904 VDD VSS sg13g2_FILL8
XSTDFILL62_1912 VDD VSS sg13g2_FILL8
XSTDFILL62_1920 VDD VSS sg13g2_FILL8
XSTDFILL62_1928 VDD VSS sg13g2_FILL8
XSTDFILL62_1936 VDD VSS sg13g2_FILL8
XSTDFILL62_1944 VDD VSS sg13g2_FILL8
XSTDFILL62_1952 VDD VSS sg13g2_FILL8
XSTDFILL62_1960 VDD VSS sg13g2_FILL8
XSTDFILL62_1968 VDD VSS sg13g2_FILL8
XSTDFILL62_1976 VDD VSS sg13g2_FILL8
XSTDFILL62_1984 VDD VSS sg13g2_FILL8
XSTDFILL62_1992 VDD VSS sg13g2_FILL8
XSTDFILL62_2000 VDD VSS sg13g2_FILL8
XSTDFILL62_2008 VDD VSS sg13g2_FILL8
XSTDFILL62_2016 VDD VSS sg13g2_FILL8
XSTDFILL62_2024 VDD VSS sg13g2_FILL8
XSTDFILL62_2032 VDD VSS sg13g2_FILL8
XSTDFILL62_2040 VDD VSS sg13g2_FILL8
XSTDFILL62_2048 VDD VSS sg13g2_FILL8
XSTDFILL62_2056 VDD VSS sg13g2_FILL8
XSTDFILL62_2064 VDD VSS sg13g2_FILL8
XSTDFILL62_2072 VDD VSS sg13g2_FILL8
XSTDFILL62_2080 VDD VSS sg13g2_FILL8
XSTDFILL62_2088 VDD VSS sg13g2_FILL8
XSTDFILL62_2096 VDD VSS sg13g2_FILL8
XSTDFILL62_2104 VDD VSS sg13g2_FILL8
XSTDFILL62_2112 VDD VSS sg13g2_FILL8
XSTDFILL62_2120 VDD VSS sg13g2_FILL8
XSTDFILL62_2128 VDD VSS sg13g2_FILL8
XSTDFILL62_2136 VDD VSS sg13g2_FILL8
XSTDFILL62_2144 VDD VSS sg13g2_FILL8
XSTDFILL62_2152 VDD VSS sg13g2_FILL8
XSTDFILL62_2160 VDD VSS sg13g2_FILL8
XSTDFILL62_2168 VDD VSS sg13g2_FILL4
XSTDFILL63_0 VDD VSS sg13g2_FILL8
XSTDFILL63_8 VDD VSS sg13g2_FILL8
XSTDFILL63_16 VDD VSS sg13g2_FILL8
XSTDFILL63_24 VDD VSS sg13g2_FILL8
XSTDFILL63_32 VDD VSS sg13g2_FILL8
XSTDFILL63_40 VDD VSS sg13g2_FILL8
XSTDFILL63_48 VDD VSS sg13g2_FILL8
XSTDFILL63_56 VDD VSS sg13g2_FILL8
XSTDFILL63_64 VDD VSS sg13g2_FILL8
XSTDFILL63_72 VDD VSS sg13g2_FILL8
XSTDFILL63_80 VDD VSS sg13g2_FILL8
XSTDFILL63_88 VDD VSS sg13g2_FILL8
XSTDFILL63_96 VDD VSS sg13g2_FILL8
XSTDFILL63_104 VDD VSS sg13g2_FILL8
XSTDFILL63_112 VDD VSS sg13g2_FILL8
XSTDFILL63_120 VDD VSS sg13g2_FILL8
XSTDFILL63_128 VDD VSS sg13g2_FILL8
XSTDFILL63_136 VDD VSS sg13g2_FILL8
XSTDFILL63_144 VDD VSS sg13g2_FILL8
XSTDFILL63_152 VDD VSS sg13g2_FILL8
XSTDFILL63_160 VDD VSS sg13g2_FILL8
XSTDFILL63_168 VDD VSS sg13g2_FILL8
XSTDFILL63_176 VDD VSS sg13g2_FILL8
XSTDFILL63_184 VDD VSS sg13g2_FILL8
XSTDFILL63_192 VDD VSS sg13g2_FILL8
XSTDFILL63_200 VDD VSS sg13g2_FILL8
XSTDFILL63_208 VDD VSS sg13g2_FILL8
XSTDFILL63_216 VDD VSS sg13g2_FILL8
XSTDFILL63_224 VDD VSS sg13g2_FILL8
XSTDFILL63_232 VDD VSS sg13g2_FILL8
XSTDFILL63_240 VDD VSS sg13g2_FILL8
XSTDFILL63_248 VDD VSS sg13g2_FILL8
XSTDFILL63_256 VDD VSS sg13g2_FILL8
XSTDFILL63_264 VDD VSS sg13g2_FILL8
XSTDFILL63_272 VDD VSS sg13g2_FILL8
XSTDFILL63_280 VDD VSS sg13g2_FILL8
XSTDFILL63_288 VDD VSS sg13g2_FILL8
XSTDFILL63_296 VDD VSS sg13g2_FILL8
XSTDFILL63_304 VDD VSS sg13g2_FILL8
XSTDFILL63_312 VDD VSS sg13g2_FILL8
XSTDFILL63_320 VDD VSS sg13g2_FILL8
XSTDFILL63_328 VDD VSS sg13g2_FILL8
XSTDFILL63_336 VDD VSS sg13g2_FILL8
XSTDFILL63_344 VDD VSS sg13g2_FILL8
XSTDFILL63_352 VDD VSS sg13g2_FILL8
XSTDFILL63_360 VDD VSS sg13g2_FILL8
XSTDFILL63_368 VDD VSS sg13g2_FILL8
XSTDFILL63_376 VDD VSS sg13g2_FILL8
XSTDFILL63_384 VDD VSS sg13g2_FILL8
XSTDFILL63_392 VDD VSS sg13g2_FILL8
XSTDFILL63_400 VDD VSS sg13g2_FILL8
XSTDFILL63_408 VDD VSS sg13g2_FILL8
XSTDFILL63_416 VDD VSS sg13g2_FILL8
XSTDFILL63_424 VDD VSS sg13g2_FILL8
XSTDFILL63_432 VDD VSS sg13g2_FILL8
XSTDFILL63_440 VDD VSS sg13g2_FILL8
XSTDFILL63_448 VDD VSS sg13g2_FILL8
XSTDFILL63_456 VDD VSS sg13g2_FILL8
XSTDFILL63_464 VDD VSS sg13g2_FILL8
XSTDFILL63_472 VDD VSS sg13g2_FILL8
XSTDFILL63_480 VDD VSS sg13g2_FILL8
XSTDFILL63_488 VDD VSS sg13g2_FILL8
XSTDFILL63_496 VDD VSS sg13g2_FILL8
XSTDFILL63_504 VDD VSS sg13g2_FILL8
XSTDFILL63_512 VDD VSS sg13g2_FILL8
XSTDFILL63_520 VDD VSS sg13g2_FILL8
XSTDFILL63_528 VDD VSS sg13g2_FILL8
XSTDFILL63_536 VDD VSS sg13g2_FILL8
XSTDFILL63_544 VDD VSS sg13g2_FILL8
XSTDFILL63_552 VDD VSS sg13g2_FILL8
XSTDFILL63_560 VDD VSS sg13g2_FILL8
XSTDFILL63_568 VDD VSS sg13g2_FILL8
XSTDFILL63_576 VDD VSS sg13g2_FILL8
XSTDFILL63_584 VDD VSS sg13g2_FILL8
XSTDFILL63_592 VDD VSS sg13g2_FILL8
XSTDFILL63_600 VDD VSS sg13g2_FILL8
XSTDFILL63_608 VDD VSS sg13g2_FILL8
XSTDFILL63_616 VDD VSS sg13g2_FILL8
XSTDFILL63_624 VDD VSS sg13g2_FILL8
XSTDFILL63_632 VDD VSS sg13g2_FILL8
XSTDFILL63_640 VDD VSS sg13g2_FILL8
XSTDFILL63_648 VDD VSS sg13g2_FILL8
XSTDFILL63_656 VDD VSS sg13g2_FILL8
XSTDFILL63_664 VDD VSS sg13g2_FILL8
XSTDFILL63_672 VDD VSS sg13g2_FILL8
XSTDFILL63_680 VDD VSS sg13g2_FILL8
XSTDFILL63_688 VDD VSS sg13g2_FILL8
XSTDFILL63_696 VDD VSS sg13g2_FILL8
XSTDFILL63_704 VDD VSS sg13g2_FILL8
XSTDFILL63_712 VDD VSS sg13g2_FILL8
XSTDFILL63_720 VDD VSS sg13g2_FILL8
XSTDFILL63_728 VDD VSS sg13g2_FILL8
XSTDFILL63_736 VDD VSS sg13g2_FILL8
XSTDFILL63_744 VDD VSS sg13g2_FILL8
XSTDFILL63_752 VDD VSS sg13g2_FILL8
XSTDFILL63_760 VDD VSS sg13g2_FILL8
XSTDFILL63_768 VDD VSS sg13g2_FILL8
XSTDFILL63_776 VDD VSS sg13g2_FILL8
XSTDFILL63_784 VDD VSS sg13g2_FILL8
XSTDFILL63_792 VDD VSS sg13g2_FILL8
XSTDFILL63_800 VDD VSS sg13g2_FILL8
XSTDFILL63_808 VDD VSS sg13g2_FILL8
XSTDFILL63_816 VDD VSS sg13g2_FILL8
XSTDFILL63_824 VDD VSS sg13g2_FILL8
XSTDFILL63_832 VDD VSS sg13g2_FILL8
XSTDFILL63_840 VDD VSS sg13g2_FILL8
XSTDFILL63_848 VDD VSS sg13g2_FILL8
XSTDFILL63_856 VDD VSS sg13g2_FILL8
XSTDFILL63_864 VDD VSS sg13g2_FILL8
XSTDFILL63_872 VDD VSS sg13g2_FILL8
XSTDFILL63_880 VDD VSS sg13g2_FILL8
XSTDFILL63_888 VDD VSS sg13g2_FILL8
XSTDFILL63_896 VDD VSS sg13g2_FILL8
XSTDFILL63_904 VDD VSS sg13g2_FILL8
XSTDFILL63_912 VDD VSS sg13g2_FILL8
XSTDFILL63_920 VDD VSS sg13g2_FILL8
XSTDFILL63_928 VDD VSS sg13g2_FILL8
XSTDFILL63_936 VDD VSS sg13g2_FILL8
XSTDFILL63_944 VDD VSS sg13g2_FILL8
XSTDFILL63_952 VDD VSS sg13g2_FILL8
XSTDFILL63_960 VDD VSS sg13g2_FILL8
XSTDFILL63_968 VDD VSS sg13g2_FILL8
XSTDFILL63_976 VDD VSS sg13g2_FILL8
XSTDFILL63_984 VDD VSS sg13g2_FILL8
XSTDFILL63_992 VDD VSS sg13g2_FILL8
XSTDFILL63_1000 VDD VSS sg13g2_FILL8
XSTDFILL63_1008 VDD VSS sg13g2_FILL8
XSTDFILL63_1016 VDD VSS sg13g2_FILL8
XSTDFILL63_1024 VDD VSS sg13g2_FILL8
XSTDFILL63_1032 VDD VSS sg13g2_FILL8
XSTDFILL63_1040 VDD VSS sg13g2_FILL8
XSTDFILL63_1048 VDD VSS sg13g2_FILL8
XSTDFILL63_1056 VDD VSS sg13g2_FILL8
XSTDFILL63_1064 VDD VSS sg13g2_FILL8
XSTDFILL63_1072 VDD VSS sg13g2_FILL8
XSTDFILL63_1080 VDD VSS sg13g2_FILL8
XSTDFILL63_1088 VDD VSS sg13g2_FILL8
XSTDFILL63_1096 VDD VSS sg13g2_FILL8
XSTDFILL63_1104 VDD VSS sg13g2_FILL8
XSTDFILL63_1112 VDD VSS sg13g2_FILL8
XSTDFILL63_1120 VDD VSS sg13g2_FILL8
XSTDFILL63_1128 VDD VSS sg13g2_FILL8
XSTDFILL63_1136 VDD VSS sg13g2_FILL8
XSTDFILL63_1144 VDD VSS sg13g2_FILL8
XSTDFILL63_1152 VDD VSS sg13g2_FILL8
XSTDFILL63_1160 VDD VSS sg13g2_FILL8
XSTDFILL63_1168 VDD VSS sg13g2_FILL8
XSTDFILL63_1176 VDD VSS sg13g2_FILL8
XSTDFILL63_1184 VDD VSS sg13g2_FILL8
XSTDFILL63_1192 VDD VSS sg13g2_FILL8
XSTDFILL63_1200 VDD VSS sg13g2_FILL8
XSTDFILL63_1208 VDD VSS sg13g2_FILL8
XSTDFILL63_1216 VDD VSS sg13g2_FILL8
XSTDFILL63_1224 VDD VSS sg13g2_FILL8
XSTDFILL63_1232 VDD VSS sg13g2_FILL8
XSTDFILL63_1240 VDD VSS sg13g2_FILL8
XSTDFILL63_1248 VDD VSS sg13g2_FILL8
XSTDFILL63_1256 VDD VSS sg13g2_FILL8
XSTDFILL63_1264 VDD VSS sg13g2_FILL8
XSTDFILL63_1272 VDD VSS sg13g2_FILL8
XSTDFILL63_1280 VDD VSS sg13g2_FILL8
XSTDFILL63_1288 VDD VSS sg13g2_FILL8
XSTDFILL63_1296 VDD VSS sg13g2_FILL8
XSTDFILL63_1304 VDD VSS sg13g2_FILL8
XSTDFILL63_1312 VDD VSS sg13g2_FILL8
XSTDFILL63_1320 VDD VSS sg13g2_FILL8
XSTDFILL63_1328 VDD VSS sg13g2_FILL8
XSTDFILL63_1336 VDD VSS sg13g2_FILL8
XSTDFILL63_1344 VDD VSS sg13g2_FILL8
XSTDFILL63_1352 VDD VSS sg13g2_FILL8
XSTDFILL63_1360 VDD VSS sg13g2_FILL8
XSTDFILL63_1368 VDD VSS sg13g2_FILL8
XSTDFILL63_1376 VDD VSS sg13g2_FILL8
XSTDFILL63_1384 VDD VSS sg13g2_FILL8
XSTDFILL63_1392 VDD VSS sg13g2_FILL8
XSTDFILL63_1400 VDD VSS sg13g2_FILL8
XSTDFILL63_1408 VDD VSS sg13g2_FILL8
XSTDFILL63_1416 VDD VSS sg13g2_FILL8
XSTDFILL63_1424 VDD VSS sg13g2_FILL8
XSTDFILL63_1432 VDD VSS sg13g2_FILL8
XSTDFILL63_1440 VDD VSS sg13g2_FILL8
XSTDFILL63_1448 VDD VSS sg13g2_FILL8
XSTDFILL63_1456 VDD VSS sg13g2_FILL8
XSTDFILL63_1464 VDD VSS sg13g2_FILL8
XSTDFILL63_1472 VDD VSS sg13g2_FILL8
XSTDFILL63_1480 VDD VSS sg13g2_FILL8
XSTDFILL63_1488 VDD VSS sg13g2_FILL8
XSTDFILL63_1496 VDD VSS sg13g2_FILL8
XSTDFILL63_1504 VDD VSS sg13g2_FILL8
XSTDFILL63_1512 VDD VSS sg13g2_FILL8
XSTDFILL63_1520 VDD VSS sg13g2_FILL8
XSTDFILL63_1528 VDD VSS sg13g2_FILL8
XSTDFILL63_1536 VDD VSS sg13g2_FILL8
XSTDFILL63_1544 VDD VSS sg13g2_FILL8
XSTDFILL63_1552 VDD VSS sg13g2_FILL8
XSTDFILL63_1560 VDD VSS sg13g2_FILL8
XSTDFILL63_1568 VDD VSS sg13g2_FILL8
XSTDFILL63_1576 VDD VSS sg13g2_FILL8
XSTDFILL63_1584 VDD VSS sg13g2_FILL8
XSTDFILL63_1592 VDD VSS sg13g2_FILL8
XSTDFILL63_1600 VDD VSS sg13g2_FILL8
XSTDFILL63_1608 VDD VSS sg13g2_FILL8
XSTDFILL63_1616 VDD VSS sg13g2_FILL8
XSTDFILL63_1624 VDD VSS sg13g2_FILL8
XSTDFILL63_1632 VDD VSS sg13g2_FILL8
XSTDFILL63_1640 VDD VSS sg13g2_FILL8
XSTDFILL63_1648 VDD VSS sg13g2_FILL8
XSTDFILL63_1656 VDD VSS sg13g2_FILL8
XSTDFILL63_1664 VDD VSS sg13g2_FILL8
XSTDFILL63_1672 VDD VSS sg13g2_FILL8
XSTDFILL63_1680 VDD VSS sg13g2_FILL8
XSTDFILL63_1688 VDD VSS sg13g2_FILL8
XSTDFILL63_1696 VDD VSS sg13g2_FILL8
XSTDFILL63_1704 VDD VSS sg13g2_FILL8
XSTDFILL63_1712 VDD VSS sg13g2_FILL8
XSTDFILL63_1720 VDD VSS sg13g2_FILL8
XSTDFILL63_1728 VDD VSS sg13g2_FILL8
XSTDFILL63_1736 VDD VSS sg13g2_FILL8
XSTDFILL63_1744 VDD VSS sg13g2_FILL8
XSTDFILL63_1752 VDD VSS sg13g2_FILL8
XSTDFILL63_1760 VDD VSS sg13g2_FILL8
XSTDFILL63_1768 VDD VSS sg13g2_FILL8
XSTDFILL63_1776 VDD VSS sg13g2_FILL8
XSTDFILL63_1784 VDD VSS sg13g2_FILL8
XSTDFILL63_1792 VDD VSS sg13g2_FILL8
XSTDFILL63_1800 VDD VSS sg13g2_FILL8
XSTDFILL63_1808 VDD VSS sg13g2_FILL8
XSTDFILL63_1816 VDD VSS sg13g2_FILL8
XSTDFILL63_1824 VDD VSS sg13g2_FILL8
XSTDFILL63_1832 VDD VSS sg13g2_FILL8
XSTDFILL63_1840 VDD VSS sg13g2_FILL8
XSTDFILL63_1848 VDD VSS sg13g2_FILL8
XSTDFILL63_1856 VDD VSS sg13g2_FILL8
XSTDFILL63_1864 VDD VSS sg13g2_FILL8
XSTDFILL63_1872 VDD VSS sg13g2_FILL8
XSTDFILL63_1880 VDD VSS sg13g2_FILL8
XSTDFILL63_1888 VDD VSS sg13g2_FILL8
XSTDFILL63_1896 VDD VSS sg13g2_FILL8
XSTDFILL63_1904 VDD VSS sg13g2_FILL8
XSTDFILL63_1912 VDD VSS sg13g2_FILL8
XSTDFILL63_1920 VDD VSS sg13g2_FILL8
XSTDFILL63_1928 VDD VSS sg13g2_FILL8
XSTDFILL63_1936 VDD VSS sg13g2_FILL8
XSTDFILL63_1944 VDD VSS sg13g2_FILL8
XSTDFILL63_1952 VDD VSS sg13g2_FILL8
XSTDFILL63_1960 VDD VSS sg13g2_FILL8
XSTDFILL63_1968 VDD VSS sg13g2_FILL8
XSTDFILL63_1976 VDD VSS sg13g2_FILL8
XSTDFILL63_1984 VDD VSS sg13g2_FILL8
XSTDFILL63_1992 VDD VSS sg13g2_FILL8
XSTDFILL63_2000 VDD VSS sg13g2_FILL8
XSTDFILL63_2008 VDD VSS sg13g2_FILL8
XSTDFILL63_2016 VDD VSS sg13g2_FILL8
XSTDFILL63_2024 VDD VSS sg13g2_FILL8
XSTDFILL63_2032 VDD VSS sg13g2_FILL8
XSTDFILL63_2040 VDD VSS sg13g2_FILL8
XSTDFILL63_2048 VDD VSS sg13g2_FILL8
XSTDFILL63_2056 VDD VSS sg13g2_FILL8
XSTDFILL63_2064 VDD VSS sg13g2_FILL8
XSTDFILL63_2072 VDD VSS sg13g2_FILL8
XSTDFILL63_2080 VDD VSS sg13g2_FILL8
XSTDFILL63_2088 VDD VSS sg13g2_FILL8
XSTDFILL63_2096 VDD VSS sg13g2_FILL8
XSTDFILL63_2104 VDD VSS sg13g2_FILL8
XSTDFILL63_2112 VDD VSS sg13g2_FILL8
XSTDFILL63_2120 VDD VSS sg13g2_FILL8
XSTDFILL63_2128 VDD VSS sg13g2_FILL8
XSTDFILL63_2136 VDD VSS sg13g2_FILL8
XSTDFILL63_2144 VDD VSS sg13g2_FILL8
XSTDFILL63_2152 VDD VSS sg13g2_FILL8
XSTDFILL63_2160 VDD VSS sg13g2_FILL8
XSTDFILL63_2168 VDD VSS sg13g2_FILL4
XSTDFILL64_0 VDD VSS sg13g2_FILL8
XSTDFILL64_8 VDD VSS sg13g2_FILL8
XSTDFILL64_16 VDD VSS sg13g2_FILL8
XSTDFILL64_24 VDD VSS sg13g2_FILL8
XSTDFILL64_32 VDD VSS sg13g2_FILL8
XSTDFILL64_40 VDD VSS sg13g2_FILL8
XSTDFILL64_48 VDD VSS sg13g2_FILL8
XSTDFILL64_56 VDD VSS sg13g2_FILL8
XSTDFILL64_64 VDD VSS sg13g2_FILL8
XSTDFILL64_72 VDD VSS sg13g2_FILL8
XSTDFILL64_80 VDD VSS sg13g2_FILL8
XSTDFILL64_88 VDD VSS sg13g2_FILL8
XSTDFILL64_96 VDD VSS sg13g2_FILL8
XSTDFILL64_104 VDD VSS sg13g2_FILL8
XSTDFILL64_112 VDD VSS sg13g2_FILL8
XSTDFILL64_120 VDD VSS sg13g2_FILL8
XSTDFILL64_128 VDD VSS sg13g2_FILL8
XSTDFILL64_136 VDD VSS sg13g2_FILL8
XSTDFILL64_144 VDD VSS sg13g2_FILL8
XSTDFILL64_152 VDD VSS sg13g2_FILL8
XSTDFILL64_160 VDD VSS sg13g2_FILL8
XSTDFILL64_168 VDD VSS sg13g2_FILL8
XSTDFILL64_176 VDD VSS sg13g2_FILL8
XSTDFILL64_184 VDD VSS sg13g2_FILL8
XSTDFILL64_192 VDD VSS sg13g2_FILL8
XSTDFILL64_200 VDD VSS sg13g2_FILL8
XSTDFILL64_208 VDD VSS sg13g2_FILL8
XSTDFILL64_216 VDD VSS sg13g2_FILL8
XSTDFILL64_224 VDD VSS sg13g2_FILL8
XSTDFILL64_232 VDD VSS sg13g2_FILL8
XSTDFILL64_240 VDD VSS sg13g2_FILL8
XSTDFILL64_248 VDD VSS sg13g2_FILL8
XSTDFILL64_256 VDD VSS sg13g2_FILL8
XSTDFILL64_264 VDD VSS sg13g2_FILL8
XSTDFILL64_272 VDD VSS sg13g2_FILL8
XSTDFILL64_280 VDD VSS sg13g2_FILL8
XSTDFILL64_288 VDD VSS sg13g2_FILL8
XSTDFILL64_296 VDD VSS sg13g2_FILL8
XSTDFILL64_304 VDD VSS sg13g2_FILL8
XSTDFILL64_312 VDD VSS sg13g2_FILL8
XSTDFILL64_320 VDD VSS sg13g2_FILL8
XSTDFILL64_328 VDD VSS sg13g2_FILL8
XSTDFILL64_336 VDD VSS sg13g2_FILL8
XSTDFILL64_344 VDD VSS sg13g2_FILL8
XSTDFILL64_352 VDD VSS sg13g2_FILL8
XSTDFILL64_360 VDD VSS sg13g2_FILL8
XSTDFILL64_368 VDD VSS sg13g2_FILL8
XSTDFILL64_376 VDD VSS sg13g2_FILL8
XSTDFILL64_384 VDD VSS sg13g2_FILL8
XSTDFILL64_392 VDD VSS sg13g2_FILL8
XSTDFILL64_400 VDD VSS sg13g2_FILL8
XSTDFILL64_408 VDD VSS sg13g2_FILL8
XSTDFILL64_416 VDD VSS sg13g2_FILL8
XSTDFILL64_424 VDD VSS sg13g2_FILL8
XSTDFILL64_432 VDD VSS sg13g2_FILL8
XSTDFILL64_440 VDD VSS sg13g2_FILL8
XSTDFILL64_448 VDD VSS sg13g2_FILL8
XSTDFILL64_456 VDD VSS sg13g2_FILL8
XSTDFILL64_464 VDD VSS sg13g2_FILL8
XSTDFILL64_472 VDD VSS sg13g2_FILL8
XSTDFILL64_480 VDD VSS sg13g2_FILL8
XSTDFILL64_488 VDD VSS sg13g2_FILL8
XSTDFILL64_496 VDD VSS sg13g2_FILL8
XSTDFILL64_504 VDD VSS sg13g2_FILL8
XSTDFILL64_512 VDD VSS sg13g2_FILL8
XSTDFILL64_520 VDD VSS sg13g2_FILL8
XSTDFILL64_528 VDD VSS sg13g2_FILL8
XSTDFILL64_536 VDD VSS sg13g2_FILL8
XSTDFILL64_544 VDD VSS sg13g2_FILL8
XSTDFILL64_552 VDD VSS sg13g2_FILL8
XSTDFILL64_560 VDD VSS sg13g2_FILL8
XSTDFILL64_568 VDD VSS sg13g2_FILL8
XSTDFILL64_576 VDD VSS sg13g2_FILL8
XSTDFILL64_584 VDD VSS sg13g2_FILL8
XSTDFILL64_592 VDD VSS sg13g2_FILL8
XSTDFILL64_600 VDD VSS sg13g2_FILL8
XSTDFILL64_608 VDD VSS sg13g2_FILL8
XSTDFILL64_616 VDD VSS sg13g2_FILL8
XSTDFILL64_624 VDD VSS sg13g2_FILL8
XSTDFILL64_632 VDD VSS sg13g2_FILL8
XSTDFILL64_640 VDD VSS sg13g2_FILL8
XSTDFILL64_648 VDD VSS sg13g2_FILL8
XSTDFILL64_656 VDD VSS sg13g2_FILL8
XSTDFILL64_664 VDD VSS sg13g2_FILL8
XSTDFILL64_672 VDD VSS sg13g2_FILL8
XSTDFILL64_680 VDD VSS sg13g2_FILL8
XSTDFILL64_688 VDD VSS sg13g2_FILL8
XSTDFILL64_696 VDD VSS sg13g2_FILL8
XSTDFILL64_704 VDD VSS sg13g2_FILL8
XSTDFILL64_712 VDD VSS sg13g2_FILL8
XSTDFILL64_720 VDD VSS sg13g2_FILL8
XSTDFILL64_728 VDD VSS sg13g2_FILL8
XSTDFILL64_736 VDD VSS sg13g2_FILL8
XSTDFILL64_744 VDD VSS sg13g2_FILL8
XSTDFILL64_752 VDD VSS sg13g2_FILL8
XSTDFILL64_760 VDD VSS sg13g2_FILL8
XSTDFILL64_768 VDD VSS sg13g2_FILL8
XSTDFILL64_776 VDD VSS sg13g2_FILL8
XSTDFILL64_784 VDD VSS sg13g2_FILL8
XSTDFILL64_792 VDD VSS sg13g2_FILL8
XSTDFILL64_800 VDD VSS sg13g2_FILL8
XSTDFILL64_808 VDD VSS sg13g2_FILL8
XSTDFILL64_816 VDD VSS sg13g2_FILL8
XSTDFILL64_824 VDD VSS sg13g2_FILL8
XSTDFILL64_832 VDD VSS sg13g2_FILL8
XSTDFILL64_840 VDD VSS sg13g2_FILL8
XSTDFILL64_848 VDD VSS sg13g2_FILL8
XSTDFILL64_856 VDD VSS sg13g2_FILL8
XSTDFILL64_864 VDD VSS sg13g2_FILL8
XSTDFILL64_872 VDD VSS sg13g2_FILL8
XSTDFILL64_880 VDD VSS sg13g2_FILL8
XSTDFILL64_888 VDD VSS sg13g2_FILL8
XSTDFILL64_896 VDD VSS sg13g2_FILL8
XSTDFILL64_904 VDD VSS sg13g2_FILL8
XSTDFILL64_912 VDD VSS sg13g2_FILL8
XSTDFILL64_920 VDD VSS sg13g2_FILL8
XSTDFILL64_928 VDD VSS sg13g2_FILL8
XSTDFILL64_936 VDD VSS sg13g2_FILL8
XSTDFILL64_944 VDD VSS sg13g2_FILL8
XSTDFILL64_952 VDD VSS sg13g2_FILL8
XSTDFILL64_960 VDD VSS sg13g2_FILL8
XSTDFILL64_968 VDD VSS sg13g2_FILL8
XSTDFILL64_976 VDD VSS sg13g2_FILL8
XSTDFILL64_984 VDD VSS sg13g2_FILL8
XSTDFILL64_992 VDD VSS sg13g2_FILL8
XSTDFILL64_1000 VDD VSS sg13g2_FILL8
XSTDFILL64_1008 VDD VSS sg13g2_FILL8
XSTDFILL64_1016 VDD VSS sg13g2_FILL8
XSTDFILL64_1024 VDD VSS sg13g2_FILL8
XSTDFILL64_1032 VDD VSS sg13g2_FILL8
XSTDFILL64_1040 VDD VSS sg13g2_FILL8
XSTDFILL64_1048 VDD VSS sg13g2_FILL8
XSTDFILL64_1056 VDD VSS sg13g2_FILL8
XSTDFILL64_1064 VDD VSS sg13g2_FILL8
XSTDFILL64_1072 VDD VSS sg13g2_FILL8
XSTDFILL64_1080 VDD VSS sg13g2_FILL8
XSTDFILL64_1088 VDD VSS sg13g2_FILL8
XSTDFILL64_1096 VDD VSS sg13g2_FILL8
XSTDFILL64_1104 VDD VSS sg13g2_FILL8
XSTDFILL64_1112 VDD VSS sg13g2_FILL8
XSTDFILL64_1120 VDD VSS sg13g2_FILL8
XSTDFILL64_1128 VDD VSS sg13g2_FILL8
XSTDFILL64_1136 VDD VSS sg13g2_FILL8
XSTDFILL64_1144 VDD VSS sg13g2_FILL8
XSTDFILL64_1152 VDD VSS sg13g2_FILL8
XSTDFILL64_1160 VDD VSS sg13g2_FILL8
XSTDFILL64_1168 VDD VSS sg13g2_FILL8
XSTDFILL64_1176 VDD VSS sg13g2_FILL8
XSTDFILL64_1184 VDD VSS sg13g2_FILL8
XSTDFILL64_1192 VDD VSS sg13g2_FILL8
XSTDFILL64_1200 VDD VSS sg13g2_FILL8
XSTDFILL64_1208 VDD VSS sg13g2_FILL8
XSTDFILL64_1216 VDD VSS sg13g2_FILL8
XSTDFILL64_1224 VDD VSS sg13g2_FILL8
XSTDFILL64_1232 VDD VSS sg13g2_FILL8
XSTDFILL64_1240 VDD VSS sg13g2_FILL8
XSTDFILL64_1248 VDD VSS sg13g2_FILL8
XSTDFILL64_1256 VDD VSS sg13g2_FILL8
XSTDFILL64_1264 VDD VSS sg13g2_FILL8
XSTDFILL64_1272 VDD VSS sg13g2_FILL8
XSTDFILL64_1280 VDD VSS sg13g2_FILL8
XSTDFILL64_1288 VDD VSS sg13g2_FILL8
XSTDFILL64_1296 VDD VSS sg13g2_FILL8
XSTDFILL64_1304 VDD VSS sg13g2_FILL8
XSTDFILL64_1312 VDD VSS sg13g2_FILL8
XSTDFILL64_1320 VDD VSS sg13g2_FILL8
XSTDFILL64_1328 VDD VSS sg13g2_FILL8
XSTDFILL64_1336 VDD VSS sg13g2_FILL8
XSTDFILL64_1344 VDD VSS sg13g2_FILL8
XSTDFILL64_1352 VDD VSS sg13g2_FILL8
XSTDFILL64_1360 VDD VSS sg13g2_FILL8
XSTDFILL64_1368 VDD VSS sg13g2_FILL8
XSTDFILL64_1376 VDD VSS sg13g2_FILL8
XSTDFILL64_1384 VDD VSS sg13g2_FILL8
XSTDFILL64_1392 VDD VSS sg13g2_FILL8
XSTDFILL64_1400 VDD VSS sg13g2_FILL8
XSTDFILL64_1408 VDD VSS sg13g2_FILL8
XSTDFILL64_1416 VDD VSS sg13g2_FILL8
XSTDFILL64_1424 VDD VSS sg13g2_FILL8
XSTDFILL64_1432 VDD VSS sg13g2_FILL8
XSTDFILL64_1440 VDD VSS sg13g2_FILL8
XSTDFILL64_1448 VDD VSS sg13g2_FILL8
XSTDFILL64_1456 VDD VSS sg13g2_FILL8
XSTDFILL64_1464 VDD VSS sg13g2_FILL8
XSTDFILL64_1472 VDD VSS sg13g2_FILL8
XSTDFILL64_1480 VDD VSS sg13g2_FILL8
XSTDFILL64_1488 VDD VSS sg13g2_FILL8
XSTDFILL64_1496 VDD VSS sg13g2_FILL8
XSTDFILL64_1504 VDD VSS sg13g2_FILL8
XSTDFILL64_1512 VDD VSS sg13g2_FILL8
XSTDFILL64_1520 VDD VSS sg13g2_FILL8
XSTDFILL64_1528 VDD VSS sg13g2_FILL8
XSTDFILL64_1536 VDD VSS sg13g2_FILL8
XSTDFILL64_1544 VDD VSS sg13g2_FILL8
XSTDFILL64_1552 VDD VSS sg13g2_FILL8
XSTDFILL64_1560 VDD VSS sg13g2_FILL8
XSTDFILL64_1568 VDD VSS sg13g2_FILL8
XSTDFILL64_1576 VDD VSS sg13g2_FILL8
XSTDFILL64_1584 VDD VSS sg13g2_FILL8
XSTDFILL64_1592 VDD VSS sg13g2_FILL8
XSTDFILL64_1600 VDD VSS sg13g2_FILL8
XSTDFILL64_1608 VDD VSS sg13g2_FILL8
XSTDFILL64_1616 VDD VSS sg13g2_FILL8
XSTDFILL64_1624 VDD VSS sg13g2_FILL8
XSTDFILL64_1632 VDD VSS sg13g2_FILL8
XSTDFILL64_1640 VDD VSS sg13g2_FILL8
XSTDFILL64_1648 VDD VSS sg13g2_FILL8
XSTDFILL64_1656 VDD VSS sg13g2_FILL8
XSTDFILL64_1664 VDD VSS sg13g2_FILL8
XSTDFILL64_1672 VDD VSS sg13g2_FILL8
XSTDFILL64_1680 VDD VSS sg13g2_FILL8
XSTDFILL64_1688 VDD VSS sg13g2_FILL8
XSTDFILL64_1696 VDD VSS sg13g2_FILL8
XSTDFILL64_1704 VDD VSS sg13g2_FILL8
XSTDFILL64_1712 VDD VSS sg13g2_FILL8
XSTDFILL64_1720 VDD VSS sg13g2_FILL8
XSTDFILL64_1728 VDD VSS sg13g2_FILL8
XSTDFILL64_1736 VDD VSS sg13g2_FILL8
XSTDFILL64_1744 VDD VSS sg13g2_FILL8
XSTDFILL64_1752 VDD VSS sg13g2_FILL8
XSTDFILL64_1760 VDD VSS sg13g2_FILL8
XSTDFILL64_1768 VDD VSS sg13g2_FILL8
XSTDFILL64_1776 VDD VSS sg13g2_FILL8
XSTDFILL64_1784 VDD VSS sg13g2_FILL8
XSTDFILL64_1792 VDD VSS sg13g2_FILL8
XSTDFILL64_1800 VDD VSS sg13g2_FILL8
XSTDFILL64_1808 VDD VSS sg13g2_FILL8
XSTDFILL64_1816 VDD VSS sg13g2_FILL8
XSTDFILL64_1824 VDD VSS sg13g2_FILL8
XSTDFILL64_1832 VDD VSS sg13g2_FILL8
XSTDFILL64_1840 VDD VSS sg13g2_FILL8
XSTDFILL64_1848 VDD VSS sg13g2_FILL8
XSTDFILL64_1856 VDD VSS sg13g2_FILL8
XSTDFILL64_1864 VDD VSS sg13g2_FILL8
XSTDFILL64_1872 VDD VSS sg13g2_FILL8
XSTDFILL64_1880 VDD VSS sg13g2_FILL8
XSTDFILL64_1888 VDD VSS sg13g2_FILL8
XSTDFILL64_1896 VDD VSS sg13g2_FILL8
XSTDFILL64_1904 VDD VSS sg13g2_FILL8
XSTDFILL64_1912 VDD VSS sg13g2_FILL8
XSTDFILL64_1920 VDD VSS sg13g2_FILL8
XSTDFILL64_1928 VDD VSS sg13g2_FILL8
XSTDFILL64_1936 VDD VSS sg13g2_FILL8
XSTDFILL64_1944 VDD VSS sg13g2_FILL8
XSTDFILL64_1952 VDD VSS sg13g2_FILL8
XSTDFILL64_1960 VDD VSS sg13g2_FILL8
XSTDFILL64_1968 VDD VSS sg13g2_FILL8
XSTDFILL64_1976 VDD VSS sg13g2_FILL8
XSTDFILL64_1984 VDD VSS sg13g2_FILL8
XSTDFILL64_1992 VDD VSS sg13g2_FILL8
XSTDFILL64_2000 VDD VSS sg13g2_FILL8
XSTDFILL64_2008 VDD VSS sg13g2_FILL8
XSTDFILL64_2016 VDD VSS sg13g2_FILL8
XSTDFILL64_2024 VDD VSS sg13g2_FILL8
XSTDFILL64_2032 VDD VSS sg13g2_FILL8
XSTDFILL64_2040 VDD VSS sg13g2_FILL8
XSTDFILL64_2048 VDD VSS sg13g2_FILL8
XSTDFILL64_2056 VDD VSS sg13g2_FILL8
XSTDFILL64_2064 VDD VSS sg13g2_FILL8
XSTDFILL64_2072 VDD VSS sg13g2_FILL8
XSTDFILL64_2080 VDD VSS sg13g2_FILL8
XSTDFILL64_2088 VDD VSS sg13g2_FILL8
XSTDFILL64_2096 VDD VSS sg13g2_FILL8
XSTDFILL64_2104 VDD VSS sg13g2_FILL8
XSTDFILL64_2112 VDD VSS sg13g2_FILL8
XSTDFILL64_2120 VDD VSS sg13g2_FILL8
XSTDFILL64_2128 VDD VSS sg13g2_FILL8
XSTDFILL64_2136 VDD VSS sg13g2_FILL8
XSTDFILL64_2144 VDD VSS sg13g2_FILL8
XSTDFILL64_2152 VDD VSS sg13g2_FILL8
XSTDFILL64_2160 VDD VSS sg13g2_FILL8
XSTDFILL64_2168 VDD VSS sg13g2_FILL4
XSTDFILL65_0 VDD VSS sg13g2_FILL8
XSTDFILL65_8 VDD VSS sg13g2_FILL8
XSTDFILL65_16 VDD VSS sg13g2_FILL8
XSTDFILL65_24 VDD VSS sg13g2_FILL8
XSTDFILL65_32 VDD VSS sg13g2_FILL8
XSTDFILL65_40 VDD VSS sg13g2_FILL8
XSTDFILL65_48 VDD VSS sg13g2_FILL8
XSTDFILL65_56 VDD VSS sg13g2_FILL8
XSTDFILL65_64 VDD VSS sg13g2_FILL8
XSTDFILL65_72 VDD VSS sg13g2_FILL8
XSTDFILL65_80 VDD VSS sg13g2_FILL8
XSTDFILL65_88 VDD VSS sg13g2_FILL8
XSTDFILL65_96 VDD VSS sg13g2_FILL8
XSTDFILL65_104 VDD VSS sg13g2_FILL8
XSTDFILL65_112 VDD VSS sg13g2_FILL8
XSTDFILL65_120 VDD VSS sg13g2_FILL8
XSTDFILL65_128 VDD VSS sg13g2_FILL8
XSTDFILL65_136 VDD VSS sg13g2_FILL8
XSTDFILL65_144 VDD VSS sg13g2_FILL8
XSTDFILL65_152 VDD VSS sg13g2_FILL8
XSTDFILL65_160 VDD VSS sg13g2_FILL8
XSTDFILL65_168 VDD VSS sg13g2_FILL8
XSTDFILL65_176 VDD VSS sg13g2_FILL8
XSTDFILL65_184 VDD VSS sg13g2_FILL8
XSTDFILL65_192 VDD VSS sg13g2_FILL8
XSTDFILL65_200 VDD VSS sg13g2_FILL8
XSTDFILL65_208 VDD VSS sg13g2_FILL8
XSTDFILL65_216 VDD VSS sg13g2_FILL8
XSTDFILL65_224 VDD VSS sg13g2_FILL8
XSTDFILL65_232 VDD VSS sg13g2_FILL8
XSTDFILL65_240 VDD VSS sg13g2_FILL8
XSTDFILL65_248 VDD VSS sg13g2_FILL8
XSTDFILL65_256 VDD VSS sg13g2_FILL8
XSTDFILL65_264 VDD VSS sg13g2_FILL8
XSTDFILL65_272 VDD VSS sg13g2_FILL8
XSTDFILL65_280 VDD VSS sg13g2_FILL8
XSTDFILL65_288 VDD VSS sg13g2_FILL8
XSTDFILL65_296 VDD VSS sg13g2_FILL8
XSTDFILL65_304 VDD VSS sg13g2_FILL8
XSTDFILL65_312 VDD VSS sg13g2_FILL8
XSTDFILL65_320 VDD VSS sg13g2_FILL8
XSTDFILL65_328 VDD VSS sg13g2_FILL8
XSTDFILL65_336 VDD VSS sg13g2_FILL8
XSTDFILL65_344 VDD VSS sg13g2_FILL8
XSTDFILL65_352 VDD VSS sg13g2_FILL8
XSTDFILL65_360 VDD VSS sg13g2_FILL8
XSTDFILL65_368 VDD VSS sg13g2_FILL8
XSTDFILL65_376 VDD VSS sg13g2_FILL8
XSTDFILL65_384 VDD VSS sg13g2_FILL8
XSTDFILL65_392 VDD VSS sg13g2_FILL8
XSTDFILL65_400 VDD VSS sg13g2_FILL8
XSTDFILL65_408 VDD VSS sg13g2_FILL8
XSTDFILL65_416 VDD VSS sg13g2_FILL8
XSTDFILL65_424 VDD VSS sg13g2_FILL8
XSTDFILL65_432 VDD VSS sg13g2_FILL8
XSTDFILL65_440 VDD VSS sg13g2_FILL8
XSTDFILL65_448 VDD VSS sg13g2_FILL8
XSTDFILL65_456 VDD VSS sg13g2_FILL8
XSTDFILL65_464 VDD VSS sg13g2_FILL8
XSTDFILL65_472 VDD VSS sg13g2_FILL8
XSTDFILL65_480 VDD VSS sg13g2_FILL8
XSTDFILL65_488 VDD VSS sg13g2_FILL8
XSTDFILL65_496 VDD VSS sg13g2_FILL8
XSTDFILL65_504 VDD VSS sg13g2_FILL8
XSTDFILL65_512 VDD VSS sg13g2_FILL8
XSTDFILL65_520 VDD VSS sg13g2_FILL8
XSTDFILL65_528 VDD VSS sg13g2_FILL8
XSTDFILL65_536 VDD VSS sg13g2_FILL8
XSTDFILL65_544 VDD VSS sg13g2_FILL8
XSTDFILL65_552 VDD VSS sg13g2_FILL8
XSTDFILL65_560 VDD VSS sg13g2_FILL8
XSTDFILL65_568 VDD VSS sg13g2_FILL8
XSTDFILL65_576 VDD VSS sg13g2_FILL8
XSTDFILL65_584 VDD VSS sg13g2_FILL8
XSTDFILL65_592 VDD VSS sg13g2_FILL8
XSTDFILL65_600 VDD VSS sg13g2_FILL8
XSTDFILL65_608 VDD VSS sg13g2_FILL8
XSTDFILL65_616 VDD VSS sg13g2_FILL8
XSTDFILL65_624 VDD VSS sg13g2_FILL8
XSTDFILL65_632 VDD VSS sg13g2_FILL8
XSTDFILL65_640 VDD VSS sg13g2_FILL8
XSTDFILL65_648 VDD VSS sg13g2_FILL8
XSTDFILL65_656 VDD VSS sg13g2_FILL8
XSTDFILL65_664 VDD VSS sg13g2_FILL8
XSTDFILL65_672 VDD VSS sg13g2_FILL8
XSTDFILL65_680 VDD VSS sg13g2_FILL8
XSTDFILL65_688 VDD VSS sg13g2_FILL8
XSTDFILL65_696 VDD VSS sg13g2_FILL8
XSTDFILL65_704 VDD VSS sg13g2_FILL8
XSTDFILL65_712 VDD VSS sg13g2_FILL8
XSTDFILL65_720 VDD VSS sg13g2_FILL8
XSTDFILL65_728 VDD VSS sg13g2_FILL8
XSTDFILL65_736 VDD VSS sg13g2_FILL8
XSTDFILL65_744 VDD VSS sg13g2_FILL8
XSTDFILL65_752 VDD VSS sg13g2_FILL8
XSTDFILL65_760 VDD VSS sg13g2_FILL8
XSTDFILL65_768 VDD VSS sg13g2_FILL8
XSTDFILL65_776 VDD VSS sg13g2_FILL8
XSTDFILL65_784 VDD VSS sg13g2_FILL8
XSTDFILL65_792 VDD VSS sg13g2_FILL8
XSTDFILL65_800 VDD VSS sg13g2_FILL8
XSTDFILL65_808 VDD VSS sg13g2_FILL8
XSTDFILL65_816 VDD VSS sg13g2_FILL8
XSTDFILL65_824 VDD VSS sg13g2_FILL8
XSTDFILL65_832 VDD VSS sg13g2_FILL8
XSTDFILL65_840 VDD VSS sg13g2_FILL8
XSTDFILL65_848 VDD VSS sg13g2_FILL8
XSTDFILL65_856 VDD VSS sg13g2_FILL8
XSTDFILL65_864 VDD VSS sg13g2_FILL8
XSTDFILL65_872 VDD VSS sg13g2_FILL8
XSTDFILL65_880 VDD VSS sg13g2_FILL8
XSTDFILL65_888 VDD VSS sg13g2_FILL8
XSTDFILL65_896 VDD VSS sg13g2_FILL8
XSTDFILL65_904 VDD VSS sg13g2_FILL8
XSTDFILL65_912 VDD VSS sg13g2_FILL8
XSTDFILL65_920 VDD VSS sg13g2_FILL8
XSTDFILL65_928 VDD VSS sg13g2_FILL8
XSTDFILL65_936 VDD VSS sg13g2_FILL8
XSTDFILL65_944 VDD VSS sg13g2_FILL8
XSTDFILL65_952 VDD VSS sg13g2_FILL8
XSTDFILL65_960 VDD VSS sg13g2_FILL8
XSTDFILL65_968 VDD VSS sg13g2_FILL8
XSTDFILL65_976 VDD VSS sg13g2_FILL8
XSTDFILL65_984 VDD VSS sg13g2_FILL8
XSTDFILL65_992 VDD VSS sg13g2_FILL8
XSTDFILL65_1000 VDD VSS sg13g2_FILL8
XSTDFILL65_1008 VDD VSS sg13g2_FILL8
XSTDFILL65_1016 VDD VSS sg13g2_FILL8
XSTDFILL65_1024 VDD VSS sg13g2_FILL8
XSTDFILL65_1032 VDD VSS sg13g2_FILL8
XSTDFILL65_1040 VDD VSS sg13g2_FILL8
XSTDFILL65_1048 VDD VSS sg13g2_FILL8
XSTDFILL65_1056 VDD VSS sg13g2_FILL8
XSTDFILL65_1064 VDD VSS sg13g2_FILL8
XSTDFILL65_1072 VDD VSS sg13g2_FILL8
XSTDFILL65_1080 VDD VSS sg13g2_FILL8
XSTDFILL65_1088 VDD VSS sg13g2_FILL8
XSTDFILL65_1096 VDD VSS sg13g2_FILL8
XSTDFILL65_1104 VDD VSS sg13g2_FILL8
XSTDFILL65_1112 VDD VSS sg13g2_FILL8
XSTDFILL65_1120 VDD VSS sg13g2_FILL8
XSTDFILL65_1128 VDD VSS sg13g2_FILL8
XSTDFILL65_1136 VDD VSS sg13g2_FILL8
XSTDFILL65_1144 VDD VSS sg13g2_FILL8
XSTDFILL65_1152 VDD VSS sg13g2_FILL8
XSTDFILL65_1160 VDD VSS sg13g2_FILL8
XSTDFILL65_1168 VDD VSS sg13g2_FILL8
XSTDFILL65_1176 VDD VSS sg13g2_FILL8
XSTDFILL65_1184 VDD VSS sg13g2_FILL8
XSTDFILL65_1192 VDD VSS sg13g2_FILL8
XSTDFILL65_1200 VDD VSS sg13g2_FILL8
XSTDFILL65_1208 VDD VSS sg13g2_FILL8
XSTDFILL65_1216 VDD VSS sg13g2_FILL8
XSTDFILL65_1224 VDD VSS sg13g2_FILL8
XSTDFILL65_1232 VDD VSS sg13g2_FILL8
XSTDFILL65_1240 VDD VSS sg13g2_FILL8
XSTDFILL65_1248 VDD VSS sg13g2_FILL8
XSTDFILL65_1256 VDD VSS sg13g2_FILL8
XSTDFILL65_1264 VDD VSS sg13g2_FILL8
XSTDFILL65_1272 VDD VSS sg13g2_FILL8
XSTDFILL65_1280 VDD VSS sg13g2_FILL8
XSTDFILL65_1288 VDD VSS sg13g2_FILL8
XSTDFILL65_1296 VDD VSS sg13g2_FILL8
XSTDFILL65_1304 VDD VSS sg13g2_FILL8
XSTDFILL65_1312 VDD VSS sg13g2_FILL8
XSTDFILL65_1320 VDD VSS sg13g2_FILL8
XSTDFILL65_1328 VDD VSS sg13g2_FILL8
XSTDFILL65_1336 VDD VSS sg13g2_FILL8
XSTDFILL65_1344 VDD VSS sg13g2_FILL8
XSTDFILL65_1352 VDD VSS sg13g2_FILL8
XSTDFILL65_1360 VDD VSS sg13g2_FILL8
XSTDFILL65_1368 VDD VSS sg13g2_FILL8
XSTDFILL65_1376 VDD VSS sg13g2_FILL8
XSTDFILL65_1384 VDD VSS sg13g2_FILL8
XSTDFILL65_1392 VDD VSS sg13g2_FILL8
XSTDFILL65_1400 VDD VSS sg13g2_FILL8
XSTDFILL65_1408 VDD VSS sg13g2_FILL8
XSTDFILL65_1416 VDD VSS sg13g2_FILL8
XSTDFILL65_1424 VDD VSS sg13g2_FILL8
XSTDFILL65_1432 VDD VSS sg13g2_FILL8
XSTDFILL65_1440 VDD VSS sg13g2_FILL8
XSTDFILL65_1448 VDD VSS sg13g2_FILL8
XSTDFILL65_1456 VDD VSS sg13g2_FILL8
XSTDFILL65_1464 VDD VSS sg13g2_FILL8
XSTDFILL65_1472 VDD VSS sg13g2_FILL8
XSTDFILL65_1480 VDD VSS sg13g2_FILL8
XSTDFILL65_1488 VDD VSS sg13g2_FILL8
XSTDFILL65_1496 VDD VSS sg13g2_FILL8
XSTDFILL65_1504 VDD VSS sg13g2_FILL8
XSTDFILL65_1512 VDD VSS sg13g2_FILL8
XSTDFILL65_1520 VDD VSS sg13g2_FILL8
XSTDFILL65_1528 VDD VSS sg13g2_FILL8
XSTDFILL65_1536 VDD VSS sg13g2_FILL8
XSTDFILL65_1544 VDD VSS sg13g2_FILL8
XSTDFILL65_1552 VDD VSS sg13g2_FILL8
XSTDFILL65_1560 VDD VSS sg13g2_FILL8
XSTDFILL65_1568 VDD VSS sg13g2_FILL8
XSTDFILL65_1576 VDD VSS sg13g2_FILL8
XSTDFILL65_1584 VDD VSS sg13g2_FILL8
XSTDFILL65_1592 VDD VSS sg13g2_FILL8
XSTDFILL65_1600 VDD VSS sg13g2_FILL8
XSTDFILL65_1608 VDD VSS sg13g2_FILL8
XSTDFILL65_1616 VDD VSS sg13g2_FILL8
XSTDFILL65_1624 VDD VSS sg13g2_FILL8
XSTDFILL65_1632 VDD VSS sg13g2_FILL8
XSTDFILL65_1640 VDD VSS sg13g2_FILL8
XSTDFILL65_1648 VDD VSS sg13g2_FILL8
XSTDFILL65_1656 VDD VSS sg13g2_FILL8
XSTDFILL65_1664 VDD VSS sg13g2_FILL8
XSTDFILL65_1672 VDD VSS sg13g2_FILL8
XSTDFILL65_1680 VDD VSS sg13g2_FILL8
XSTDFILL65_1688 VDD VSS sg13g2_FILL8
XSTDFILL65_1696 VDD VSS sg13g2_FILL8
XSTDFILL65_1704 VDD VSS sg13g2_FILL8
XSTDFILL65_1712 VDD VSS sg13g2_FILL8
XSTDFILL65_1720 VDD VSS sg13g2_FILL8
XSTDFILL65_1728 VDD VSS sg13g2_FILL8
XSTDFILL65_1736 VDD VSS sg13g2_FILL8
XSTDFILL65_1744 VDD VSS sg13g2_FILL8
XSTDFILL65_1752 VDD VSS sg13g2_FILL8
XSTDFILL65_1760 VDD VSS sg13g2_FILL8
XSTDFILL65_1768 VDD VSS sg13g2_FILL8
XSTDFILL65_1776 VDD VSS sg13g2_FILL8
XSTDFILL65_1784 VDD VSS sg13g2_FILL8
XSTDFILL65_1792 VDD VSS sg13g2_FILL8
XSTDFILL65_1800 VDD VSS sg13g2_FILL8
XSTDFILL65_1808 VDD VSS sg13g2_FILL8
XSTDFILL65_1816 VDD VSS sg13g2_FILL8
XSTDFILL65_1824 VDD VSS sg13g2_FILL8
XSTDFILL65_1832 VDD VSS sg13g2_FILL8
XSTDFILL65_1840 VDD VSS sg13g2_FILL8
XSTDFILL65_1848 VDD VSS sg13g2_FILL8
XSTDFILL65_1856 VDD VSS sg13g2_FILL8
XSTDFILL65_1864 VDD VSS sg13g2_FILL8
XSTDFILL65_1872 VDD VSS sg13g2_FILL8
XSTDFILL65_1880 VDD VSS sg13g2_FILL8
XSTDFILL65_1888 VDD VSS sg13g2_FILL8
XSTDFILL65_1896 VDD VSS sg13g2_FILL8
XSTDFILL65_1904 VDD VSS sg13g2_FILL8
XSTDFILL65_1912 VDD VSS sg13g2_FILL8
XSTDFILL65_1920 VDD VSS sg13g2_FILL8
XSTDFILL65_1928 VDD VSS sg13g2_FILL8
XSTDFILL65_1936 VDD VSS sg13g2_FILL8
XSTDFILL65_1944 VDD VSS sg13g2_FILL8
XSTDFILL65_1952 VDD VSS sg13g2_FILL8
XSTDFILL65_1960 VDD VSS sg13g2_FILL8
XSTDFILL65_1968 VDD VSS sg13g2_FILL8
XSTDFILL65_1976 VDD VSS sg13g2_FILL8
XSTDFILL65_1984 VDD VSS sg13g2_FILL8
XSTDFILL65_1992 VDD VSS sg13g2_FILL8
XSTDFILL65_2000 VDD VSS sg13g2_FILL8
XSTDFILL65_2008 VDD VSS sg13g2_FILL8
XSTDFILL65_2016 VDD VSS sg13g2_FILL8
XSTDFILL65_2024 VDD VSS sg13g2_FILL8
XSTDFILL65_2032 VDD VSS sg13g2_FILL8
XSTDFILL65_2040 VDD VSS sg13g2_FILL8
XSTDFILL65_2048 VDD VSS sg13g2_FILL8
XSTDFILL65_2056 VDD VSS sg13g2_FILL8
XSTDFILL65_2064 VDD VSS sg13g2_FILL8
XSTDFILL65_2072 VDD VSS sg13g2_FILL8
XSTDFILL65_2080 VDD VSS sg13g2_FILL8
XSTDFILL65_2088 VDD VSS sg13g2_FILL8
XSTDFILL65_2096 VDD VSS sg13g2_FILL8
XSTDFILL65_2104 VDD VSS sg13g2_FILL8
XSTDFILL65_2112 VDD VSS sg13g2_FILL8
XSTDFILL65_2120 VDD VSS sg13g2_FILL8
XSTDFILL65_2128 VDD VSS sg13g2_FILL8
XSTDFILL65_2136 VDD VSS sg13g2_FILL8
XSTDFILL65_2144 VDD VSS sg13g2_FILL8
XSTDFILL65_2152 VDD VSS sg13g2_FILL8
XSTDFILL65_2160 VDD VSS sg13g2_FILL8
XSTDFILL65_2168 VDD VSS sg13g2_FILL4
XSTDFILL66_0 VDD VSS sg13g2_FILL8
XSTDFILL66_8 VDD VSS sg13g2_FILL8
XSTDFILL66_16 VDD VSS sg13g2_FILL8
XSTDFILL66_24 VDD VSS sg13g2_FILL8
XSTDFILL66_32 VDD VSS sg13g2_FILL8
XSTDFILL66_40 VDD VSS sg13g2_FILL8
XSTDFILL66_48 VDD VSS sg13g2_FILL8
XSTDFILL66_56 VDD VSS sg13g2_FILL8
XSTDFILL66_64 VDD VSS sg13g2_FILL8
XSTDFILL66_72 VDD VSS sg13g2_FILL8
XSTDFILL66_80 VDD VSS sg13g2_FILL8
XSTDFILL66_88 VDD VSS sg13g2_FILL8
XSTDFILL66_96 VDD VSS sg13g2_FILL8
XSTDFILL66_104 VDD VSS sg13g2_FILL8
XSTDFILL66_112 VDD VSS sg13g2_FILL8
XSTDFILL66_120 VDD VSS sg13g2_FILL8
XSTDFILL66_128 VDD VSS sg13g2_FILL8
XSTDFILL66_136 VDD VSS sg13g2_FILL8
XSTDFILL66_144 VDD VSS sg13g2_FILL8
XSTDFILL66_152 VDD VSS sg13g2_FILL8
XSTDFILL66_160 VDD VSS sg13g2_FILL8
XSTDFILL66_168 VDD VSS sg13g2_FILL8
XSTDFILL66_176 VDD VSS sg13g2_FILL8
XSTDFILL66_184 VDD VSS sg13g2_FILL8
XSTDFILL66_192 VDD VSS sg13g2_FILL8
XSTDFILL66_200 VDD VSS sg13g2_FILL8
XSTDFILL66_208 VDD VSS sg13g2_FILL8
XSTDFILL66_216 VDD VSS sg13g2_FILL8
XSTDFILL66_224 VDD VSS sg13g2_FILL8
XSTDFILL66_232 VDD VSS sg13g2_FILL8
XSTDFILL66_240 VDD VSS sg13g2_FILL8
XSTDFILL66_248 VDD VSS sg13g2_FILL8
XSTDFILL66_256 VDD VSS sg13g2_FILL8
XSTDFILL66_264 VDD VSS sg13g2_FILL8
XSTDFILL66_272 VDD VSS sg13g2_FILL8
XSTDFILL66_280 VDD VSS sg13g2_FILL8
XSTDFILL66_288 VDD VSS sg13g2_FILL8
XSTDFILL66_296 VDD VSS sg13g2_FILL8
XSTDFILL66_304 VDD VSS sg13g2_FILL8
XSTDFILL66_312 VDD VSS sg13g2_FILL8
XSTDFILL66_320 VDD VSS sg13g2_FILL8
XSTDFILL66_328 VDD VSS sg13g2_FILL8
XSTDFILL66_336 VDD VSS sg13g2_FILL8
XSTDFILL66_344 VDD VSS sg13g2_FILL8
XSTDFILL66_352 VDD VSS sg13g2_FILL8
XSTDFILL66_360 VDD VSS sg13g2_FILL8
XSTDFILL66_368 VDD VSS sg13g2_FILL8
XSTDFILL66_376 VDD VSS sg13g2_FILL8
XSTDFILL66_384 VDD VSS sg13g2_FILL8
XSTDFILL66_392 VDD VSS sg13g2_FILL8
XSTDFILL66_400 VDD VSS sg13g2_FILL8
XSTDFILL66_408 VDD VSS sg13g2_FILL8
XSTDFILL66_416 VDD VSS sg13g2_FILL8
XSTDFILL66_424 VDD VSS sg13g2_FILL8
XSTDFILL66_432 VDD VSS sg13g2_FILL8
XSTDFILL66_440 VDD VSS sg13g2_FILL8
XSTDFILL66_448 VDD VSS sg13g2_FILL8
XSTDFILL66_456 VDD VSS sg13g2_FILL8
XSTDFILL66_464 VDD VSS sg13g2_FILL8
XSTDFILL66_472 VDD VSS sg13g2_FILL8
XSTDFILL66_480 VDD VSS sg13g2_FILL8
XSTDFILL66_488 VDD VSS sg13g2_FILL8
XSTDFILL66_496 VDD VSS sg13g2_FILL8
XSTDFILL66_504 VDD VSS sg13g2_FILL8
XSTDFILL66_512 VDD VSS sg13g2_FILL8
XSTDFILL66_520 VDD VSS sg13g2_FILL8
XSTDFILL66_528 VDD VSS sg13g2_FILL8
XSTDFILL66_536 VDD VSS sg13g2_FILL8
XSTDFILL66_544 VDD VSS sg13g2_FILL8
XSTDFILL66_552 VDD VSS sg13g2_FILL8
XSTDFILL66_560 VDD VSS sg13g2_FILL8
XSTDFILL66_568 VDD VSS sg13g2_FILL8
XSTDFILL66_576 VDD VSS sg13g2_FILL8
XSTDFILL66_584 VDD VSS sg13g2_FILL8
XSTDFILL66_592 VDD VSS sg13g2_FILL8
XSTDFILL66_600 VDD VSS sg13g2_FILL8
XSTDFILL66_608 VDD VSS sg13g2_FILL8
XSTDFILL66_616 VDD VSS sg13g2_FILL8
XSTDFILL66_624 VDD VSS sg13g2_FILL8
XSTDFILL66_632 VDD VSS sg13g2_FILL8
XSTDFILL66_640 VDD VSS sg13g2_FILL8
XSTDFILL66_648 VDD VSS sg13g2_FILL8
XSTDFILL66_656 VDD VSS sg13g2_FILL8
XSTDFILL66_664 VDD VSS sg13g2_FILL8
XSTDFILL66_672 VDD VSS sg13g2_FILL8
XSTDFILL66_680 VDD VSS sg13g2_FILL8
XSTDFILL66_688 VDD VSS sg13g2_FILL8
XSTDFILL66_696 VDD VSS sg13g2_FILL8
XSTDFILL66_704 VDD VSS sg13g2_FILL8
XSTDFILL66_712 VDD VSS sg13g2_FILL8
XSTDFILL66_720 VDD VSS sg13g2_FILL8
XSTDFILL66_728 VDD VSS sg13g2_FILL8
XSTDFILL66_736 VDD VSS sg13g2_FILL8
XSTDFILL66_744 VDD VSS sg13g2_FILL8
XSTDFILL66_752 VDD VSS sg13g2_FILL8
XSTDFILL66_760 VDD VSS sg13g2_FILL8
XSTDFILL66_768 VDD VSS sg13g2_FILL8
XSTDFILL66_776 VDD VSS sg13g2_FILL8
XSTDFILL66_784 VDD VSS sg13g2_FILL8
XSTDFILL66_792 VDD VSS sg13g2_FILL8
XSTDFILL66_800 VDD VSS sg13g2_FILL8
XSTDFILL66_808 VDD VSS sg13g2_FILL8
XSTDFILL66_816 VDD VSS sg13g2_FILL8
XSTDFILL66_824 VDD VSS sg13g2_FILL8
XSTDFILL66_832 VDD VSS sg13g2_FILL8
XSTDFILL66_840 VDD VSS sg13g2_FILL8
XSTDFILL66_848 VDD VSS sg13g2_FILL8
XSTDFILL66_856 VDD VSS sg13g2_FILL8
XSTDFILL66_864 VDD VSS sg13g2_FILL8
XSTDFILL66_872 VDD VSS sg13g2_FILL8
XSTDFILL66_880 VDD VSS sg13g2_FILL8
XSTDFILL66_888 VDD VSS sg13g2_FILL8
XSTDFILL66_896 VDD VSS sg13g2_FILL8
XSTDFILL66_904 VDD VSS sg13g2_FILL8
XSTDFILL66_912 VDD VSS sg13g2_FILL8
XSTDFILL66_920 VDD VSS sg13g2_FILL8
XSTDFILL66_928 VDD VSS sg13g2_FILL8
XSTDFILL66_936 VDD VSS sg13g2_FILL8
XSTDFILL66_944 VDD VSS sg13g2_FILL8
XSTDFILL66_952 VDD VSS sg13g2_FILL8
XSTDFILL66_960 VDD VSS sg13g2_FILL8
XSTDFILL66_968 VDD VSS sg13g2_FILL8
XSTDFILL66_976 VDD VSS sg13g2_FILL8
XSTDFILL66_984 VDD VSS sg13g2_FILL8
XSTDFILL66_992 VDD VSS sg13g2_FILL8
XSTDFILL66_1000 VDD VSS sg13g2_FILL8
XSTDFILL66_1008 VDD VSS sg13g2_FILL8
XSTDFILL66_1016 VDD VSS sg13g2_FILL8
XSTDFILL66_1024 VDD VSS sg13g2_FILL8
XSTDFILL66_1032 VDD VSS sg13g2_FILL8
XSTDFILL66_1040 VDD VSS sg13g2_FILL8
XSTDFILL66_1048 VDD VSS sg13g2_FILL8
XSTDFILL66_1056 VDD VSS sg13g2_FILL8
XSTDFILL66_1064 VDD VSS sg13g2_FILL8
XSTDFILL66_1072 VDD VSS sg13g2_FILL8
XSTDFILL66_1080 VDD VSS sg13g2_FILL8
XSTDFILL66_1088 VDD VSS sg13g2_FILL8
XSTDFILL66_1096 VDD VSS sg13g2_FILL8
XSTDFILL66_1104 VDD VSS sg13g2_FILL8
XSTDFILL66_1112 VDD VSS sg13g2_FILL8
XSTDFILL66_1120 VDD VSS sg13g2_FILL8
XSTDFILL66_1128 VDD VSS sg13g2_FILL8
XSTDFILL66_1136 VDD VSS sg13g2_FILL8
XSTDFILL66_1144 VDD VSS sg13g2_FILL8
XSTDFILL66_1152 VDD VSS sg13g2_FILL8
XSTDFILL66_1160 VDD VSS sg13g2_FILL8
XSTDFILL66_1168 VDD VSS sg13g2_FILL8
XSTDFILL66_1176 VDD VSS sg13g2_FILL8
XSTDFILL66_1184 VDD VSS sg13g2_FILL8
XSTDFILL66_1192 VDD VSS sg13g2_FILL8
XSTDFILL66_1200 VDD VSS sg13g2_FILL8
XSTDFILL66_1208 VDD VSS sg13g2_FILL8
XSTDFILL66_1216 VDD VSS sg13g2_FILL8
XSTDFILL66_1224 VDD VSS sg13g2_FILL8
XSTDFILL66_1232 VDD VSS sg13g2_FILL8
XSTDFILL66_1240 VDD VSS sg13g2_FILL8
XSTDFILL66_1248 VDD VSS sg13g2_FILL8
XSTDFILL66_1256 VDD VSS sg13g2_FILL8
XSTDFILL66_1264 VDD VSS sg13g2_FILL8
XSTDFILL66_1272 VDD VSS sg13g2_FILL8
XSTDFILL66_1280 VDD VSS sg13g2_FILL8
XSTDFILL66_1288 VDD VSS sg13g2_FILL8
XSTDFILL66_1296 VDD VSS sg13g2_FILL8
XSTDFILL66_1304 VDD VSS sg13g2_FILL8
XSTDFILL66_1312 VDD VSS sg13g2_FILL8
XSTDFILL66_1320 VDD VSS sg13g2_FILL8
XSTDFILL66_1328 VDD VSS sg13g2_FILL8
XSTDFILL66_1336 VDD VSS sg13g2_FILL8
XSTDFILL66_1344 VDD VSS sg13g2_FILL8
XSTDFILL66_1352 VDD VSS sg13g2_FILL8
XSTDFILL66_1360 VDD VSS sg13g2_FILL8
XSTDFILL66_1368 VDD VSS sg13g2_FILL8
XSTDFILL66_1376 VDD VSS sg13g2_FILL8
XSTDFILL66_1384 VDD VSS sg13g2_FILL8
XSTDFILL66_1392 VDD VSS sg13g2_FILL8
XSTDFILL66_1400 VDD VSS sg13g2_FILL8
XSTDFILL66_1408 VDD VSS sg13g2_FILL8
XSTDFILL66_1416 VDD VSS sg13g2_FILL8
XSTDFILL66_1424 VDD VSS sg13g2_FILL8
XSTDFILL66_1432 VDD VSS sg13g2_FILL8
XSTDFILL66_1440 VDD VSS sg13g2_FILL8
XSTDFILL66_1448 VDD VSS sg13g2_FILL8
XSTDFILL66_1456 VDD VSS sg13g2_FILL8
XSTDFILL66_1464 VDD VSS sg13g2_FILL8
XSTDFILL66_1472 VDD VSS sg13g2_FILL8
XSTDFILL66_1480 VDD VSS sg13g2_FILL8
XSTDFILL66_1488 VDD VSS sg13g2_FILL8
XSTDFILL66_1496 VDD VSS sg13g2_FILL8
XSTDFILL66_1504 VDD VSS sg13g2_FILL8
XSTDFILL66_1512 VDD VSS sg13g2_FILL8
XSTDFILL66_1520 VDD VSS sg13g2_FILL8
XSTDFILL66_1528 VDD VSS sg13g2_FILL8
XSTDFILL66_1536 VDD VSS sg13g2_FILL8
XSTDFILL66_1544 VDD VSS sg13g2_FILL8
XSTDFILL66_1552 VDD VSS sg13g2_FILL8
XSTDFILL66_1560 VDD VSS sg13g2_FILL8
XSTDFILL66_1568 VDD VSS sg13g2_FILL8
XSTDFILL66_1576 VDD VSS sg13g2_FILL8
XSTDFILL66_1584 VDD VSS sg13g2_FILL8
XSTDFILL66_1592 VDD VSS sg13g2_FILL8
XSTDFILL66_1600 VDD VSS sg13g2_FILL8
XSTDFILL66_1608 VDD VSS sg13g2_FILL8
XSTDFILL66_1616 VDD VSS sg13g2_FILL8
XSTDFILL66_1624 VDD VSS sg13g2_FILL8
XSTDFILL66_1632 VDD VSS sg13g2_FILL8
XSTDFILL66_1640 VDD VSS sg13g2_FILL8
XSTDFILL66_1648 VDD VSS sg13g2_FILL8
XSTDFILL66_1656 VDD VSS sg13g2_FILL8
XSTDFILL66_1664 VDD VSS sg13g2_FILL8
XSTDFILL66_1672 VDD VSS sg13g2_FILL8
XSTDFILL66_1680 VDD VSS sg13g2_FILL8
XSTDFILL66_1688 VDD VSS sg13g2_FILL8
XSTDFILL66_1696 VDD VSS sg13g2_FILL8
XSTDFILL66_1704 VDD VSS sg13g2_FILL8
XSTDFILL66_1712 VDD VSS sg13g2_FILL8
XSTDFILL66_1720 VDD VSS sg13g2_FILL8
XSTDFILL66_1728 VDD VSS sg13g2_FILL8
XSTDFILL66_1736 VDD VSS sg13g2_FILL8
XSTDFILL66_1744 VDD VSS sg13g2_FILL8
XSTDFILL66_1752 VDD VSS sg13g2_FILL8
XSTDFILL66_1760 VDD VSS sg13g2_FILL8
XSTDFILL66_1768 VDD VSS sg13g2_FILL8
XSTDFILL66_1776 VDD VSS sg13g2_FILL8
XSTDFILL66_1784 VDD VSS sg13g2_FILL8
XSTDFILL66_1792 VDD VSS sg13g2_FILL8
XSTDFILL66_1800 VDD VSS sg13g2_FILL8
XSTDFILL66_1808 VDD VSS sg13g2_FILL8
XSTDFILL66_1816 VDD VSS sg13g2_FILL8
XSTDFILL66_1824 VDD VSS sg13g2_FILL8
XSTDFILL66_1832 VDD VSS sg13g2_FILL8
XSTDFILL66_1840 VDD VSS sg13g2_FILL8
XSTDFILL66_1848 VDD VSS sg13g2_FILL8
XSTDFILL66_1856 VDD VSS sg13g2_FILL8
XSTDFILL66_1864 VDD VSS sg13g2_FILL8
XSTDFILL66_1872 VDD VSS sg13g2_FILL8
XSTDFILL66_1880 VDD VSS sg13g2_FILL8
XSTDFILL66_1888 VDD VSS sg13g2_FILL8
XSTDFILL66_1896 VDD VSS sg13g2_FILL8
XSTDFILL66_1904 VDD VSS sg13g2_FILL8
XSTDFILL66_1912 VDD VSS sg13g2_FILL8
XSTDFILL66_1920 VDD VSS sg13g2_FILL8
XSTDFILL66_1928 VDD VSS sg13g2_FILL8
XSTDFILL66_1936 VDD VSS sg13g2_FILL8
XSTDFILL66_1944 VDD VSS sg13g2_FILL8
XSTDFILL66_1952 VDD VSS sg13g2_FILL8
XSTDFILL66_1960 VDD VSS sg13g2_FILL8
XSTDFILL66_1968 VDD VSS sg13g2_FILL8
XSTDFILL66_1976 VDD VSS sg13g2_FILL8
XSTDFILL66_1984 VDD VSS sg13g2_FILL8
XSTDFILL66_1992 VDD VSS sg13g2_FILL8
XSTDFILL66_2000 VDD VSS sg13g2_FILL8
XSTDFILL66_2008 VDD VSS sg13g2_FILL8
XSTDFILL66_2016 VDD VSS sg13g2_FILL8
XSTDFILL66_2024 VDD VSS sg13g2_FILL8
XSTDFILL66_2032 VDD VSS sg13g2_FILL8
XSTDFILL66_2040 VDD VSS sg13g2_FILL8
XSTDFILL66_2048 VDD VSS sg13g2_FILL8
XSTDFILL66_2056 VDD VSS sg13g2_FILL8
XSTDFILL66_2064 VDD VSS sg13g2_FILL8
XSTDFILL66_2072 VDD VSS sg13g2_FILL8
XSTDFILL66_2080 VDD VSS sg13g2_FILL8
XSTDFILL66_2088 VDD VSS sg13g2_FILL8
XSTDFILL66_2096 VDD VSS sg13g2_FILL8
XSTDFILL66_2104 VDD VSS sg13g2_FILL8
XSTDFILL66_2112 VDD VSS sg13g2_FILL8
XSTDFILL66_2120 VDD VSS sg13g2_FILL8
XSTDFILL66_2128 VDD VSS sg13g2_FILL8
XSTDFILL66_2136 VDD VSS sg13g2_FILL8
XSTDFILL66_2144 VDD VSS sg13g2_FILL8
XSTDFILL66_2152 VDD VSS sg13g2_FILL8
XSTDFILL66_2160 VDD VSS sg13g2_FILL8
XSTDFILL66_2168 VDD VSS sg13g2_FILL4
XSTDFILL67_0 VDD VSS sg13g2_FILL8
XSTDFILL67_8 VDD VSS sg13g2_FILL8
XSTDFILL67_16 VDD VSS sg13g2_FILL8
XSTDFILL67_24 VDD VSS sg13g2_FILL8
XSTDFILL67_32 VDD VSS sg13g2_FILL8
XSTDFILL67_40 VDD VSS sg13g2_FILL8
XSTDFILL67_48 VDD VSS sg13g2_FILL8
XSTDFILL67_56 VDD VSS sg13g2_FILL8
XSTDFILL67_64 VDD VSS sg13g2_FILL8
XSTDFILL67_72 VDD VSS sg13g2_FILL8
XSTDFILL67_80 VDD VSS sg13g2_FILL8
XSTDFILL67_88 VDD VSS sg13g2_FILL8
XSTDFILL67_96 VDD VSS sg13g2_FILL8
XSTDFILL67_104 VDD VSS sg13g2_FILL8
XSTDFILL67_112 VDD VSS sg13g2_FILL8
XSTDFILL67_120 VDD VSS sg13g2_FILL8
XSTDFILL67_128 VDD VSS sg13g2_FILL8
XSTDFILL67_136 VDD VSS sg13g2_FILL8
XSTDFILL67_144 VDD VSS sg13g2_FILL8
XSTDFILL67_152 VDD VSS sg13g2_FILL8
XSTDFILL67_160 VDD VSS sg13g2_FILL8
XSTDFILL67_168 VDD VSS sg13g2_FILL8
XSTDFILL67_176 VDD VSS sg13g2_FILL8
XSTDFILL67_184 VDD VSS sg13g2_FILL8
XSTDFILL67_192 VDD VSS sg13g2_FILL8
XSTDFILL67_200 VDD VSS sg13g2_FILL8
XSTDFILL67_208 VDD VSS sg13g2_FILL8
XSTDFILL67_216 VDD VSS sg13g2_FILL8
XSTDFILL67_224 VDD VSS sg13g2_FILL8
XSTDFILL67_232 VDD VSS sg13g2_FILL8
XSTDFILL67_240 VDD VSS sg13g2_FILL8
XSTDFILL67_248 VDD VSS sg13g2_FILL8
XSTDFILL67_256 VDD VSS sg13g2_FILL8
XSTDFILL67_264 VDD VSS sg13g2_FILL8
XSTDFILL67_272 VDD VSS sg13g2_FILL8
XSTDFILL67_280 VDD VSS sg13g2_FILL8
XSTDFILL67_288 VDD VSS sg13g2_FILL8
XSTDFILL67_296 VDD VSS sg13g2_FILL8
XSTDFILL67_304 VDD VSS sg13g2_FILL8
XSTDFILL67_312 VDD VSS sg13g2_FILL8
XSTDFILL67_320 VDD VSS sg13g2_FILL8
XSTDFILL67_328 VDD VSS sg13g2_FILL8
XSTDFILL67_336 VDD VSS sg13g2_FILL8
XSTDFILL67_344 VDD VSS sg13g2_FILL8
XSTDFILL67_352 VDD VSS sg13g2_FILL8
XSTDFILL67_360 VDD VSS sg13g2_FILL8
XSTDFILL67_368 VDD VSS sg13g2_FILL8
XSTDFILL67_376 VDD VSS sg13g2_FILL8
XSTDFILL67_384 VDD VSS sg13g2_FILL8
XSTDFILL67_392 VDD VSS sg13g2_FILL8
XSTDFILL67_400 VDD VSS sg13g2_FILL8
XSTDFILL67_408 VDD VSS sg13g2_FILL8
XSTDFILL67_416 VDD VSS sg13g2_FILL8
XSTDFILL67_424 VDD VSS sg13g2_FILL8
XSTDFILL67_432 VDD VSS sg13g2_FILL8
XSTDFILL67_440 VDD VSS sg13g2_FILL8
XSTDFILL67_448 VDD VSS sg13g2_FILL8
XSTDFILL67_456 VDD VSS sg13g2_FILL8
XSTDFILL67_464 VDD VSS sg13g2_FILL8
XSTDFILL67_472 VDD VSS sg13g2_FILL8
XSTDFILL67_480 VDD VSS sg13g2_FILL8
XSTDFILL67_488 VDD VSS sg13g2_FILL8
XSTDFILL67_496 VDD VSS sg13g2_FILL8
XSTDFILL67_504 VDD VSS sg13g2_FILL8
XSTDFILL67_512 VDD VSS sg13g2_FILL8
XSTDFILL67_520 VDD VSS sg13g2_FILL8
XSTDFILL67_528 VDD VSS sg13g2_FILL8
XSTDFILL67_536 VDD VSS sg13g2_FILL8
XSTDFILL67_544 VDD VSS sg13g2_FILL8
XSTDFILL67_552 VDD VSS sg13g2_FILL8
XSTDFILL67_560 VDD VSS sg13g2_FILL8
XSTDFILL67_568 VDD VSS sg13g2_FILL8
XSTDFILL67_576 VDD VSS sg13g2_FILL8
XSTDFILL67_584 VDD VSS sg13g2_FILL8
XSTDFILL67_592 VDD VSS sg13g2_FILL8
XSTDFILL67_600 VDD VSS sg13g2_FILL8
XSTDFILL67_608 VDD VSS sg13g2_FILL8
XSTDFILL67_616 VDD VSS sg13g2_FILL8
XSTDFILL67_624 VDD VSS sg13g2_FILL8
XSTDFILL67_632 VDD VSS sg13g2_FILL8
XSTDFILL67_640 VDD VSS sg13g2_FILL8
XSTDFILL67_648 VDD VSS sg13g2_FILL8
XSTDFILL67_656 VDD VSS sg13g2_FILL8
XSTDFILL67_664 VDD VSS sg13g2_FILL8
XSTDFILL67_672 VDD VSS sg13g2_FILL8
XSTDFILL67_680 VDD VSS sg13g2_FILL8
XSTDFILL67_688 VDD VSS sg13g2_FILL8
XSTDFILL67_696 VDD VSS sg13g2_FILL8
XSTDFILL67_704 VDD VSS sg13g2_FILL8
XSTDFILL67_712 VDD VSS sg13g2_FILL8
XSTDFILL67_720 VDD VSS sg13g2_FILL8
XSTDFILL67_728 VDD VSS sg13g2_FILL8
XSTDFILL67_736 VDD VSS sg13g2_FILL8
XSTDFILL67_744 VDD VSS sg13g2_FILL8
XSTDFILL67_752 VDD VSS sg13g2_FILL8
XSTDFILL67_760 VDD VSS sg13g2_FILL8
XSTDFILL67_768 VDD VSS sg13g2_FILL8
XSTDFILL67_776 VDD VSS sg13g2_FILL8
XSTDFILL67_784 VDD VSS sg13g2_FILL8
XSTDFILL67_792 VDD VSS sg13g2_FILL8
XSTDFILL67_800 VDD VSS sg13g2_FILL8
XSTDFILL67_808 VDD VSS sg13g2_FILL8
XSTDFILL67_816 VDD VSS sg13g2_FILL8
XSTDFILL67_824 VDD VSS sg13g2_FILL8
XSTDFILL67_832 VDD VSS sg13g2_FILL8
XSTDFILL67_840 VDD VSS sg13g2_FILL8
XSTDFILL67_848 VDD VSS sg13g2_FILL8
XSTDFILL67_856 VDD VSS sg13g2_FILL8
XSTDFILL67_864 VDD VSS sg13g2_FILL8
XSTDFILL67_872 VDD VSS sg13g2_FILL8
XSTDFILL67_880 VDD VSS sg13g2_FILL8
XSTDFILL67_888 VDD VSS sg13g2_FILL8
XSTDFILL67_896 VDD VSS sg13g2_FILL8
XSTDFILL67_904 VDD VSS sg13g2_FILL8
XSTDFILL67_912 VDD VSS sg13g2_FILL8
XSTDFILL67_920 VDD VSS sg13g2_FILL8
XSTDFILL67_928 VDD VSS sg13g2_FILL8
XSTDFILL67_936 VDD VSS sg13g2_FILL8
XSTDFILL67_944 VDD VSS sg13g2_FILL8
XSTDFILL67_952 VDD VSS sg13g2_FILL8
XSTDFILL67_960 VDD VSS sg13g2_FILL8
XSTDFILL67_968 VDD VSS sg13g2_FILL8
XSTDFILL67_976 VDD VSS sg13g2_FILL8
XSTDFILL67_984 VDD VSS sg13g2_FILL8
XSTDFILL67_992 VDD VSS sg13g2_FILL8
XSTDFILL67_1000 VDD VSS sg13g2_FILL8
XSTDFILL67_1008 VDD VSS sg13g2_FILL8
XSTDFILL67_1016 VDD VSS sg13g2_FILL8
XSTDFILL67_1024 VDD VSS sg13g2_FILL8
XSTDFILL67_1032 VDD VSS sg13g2_FILL8
XSTDFILL67_1040 VDD VSS sg13g2_FILL8
XSTDFILL67_1048 VDD VSS sg13g2_FILL8
XSTDFILL67_1056 VDD VSS sg13g2_FILL8
XSTDFILL67_1064 VDD VSS sg13g2_FILL8
XSTDFILL67_1072 VDD VSS sg13g2_FILL8
XSTDFILL67_1080 VDD VSS sg13g2_FILL8
XSTDFILL67_1088 VDD VSS sg13g2_FILL8
XSTDFILL67_1096 VDD VSS sg13g2_FILL8
XSTDFILL67_1104 VDD VSS sg13g2_FILL8
XSTDFILL67_1112 VDD VSS sg13g2_FILL8
XSTDFILL67_1120 VDD VSS sg13g2_FILL8
XSTDFILL67_1128 VDD VSS sg13g2_FILL8
XSTDFILL67_1136 VDD VSS sg13g2_FILL8
XSTDFILL67_1144 VDD VSS sg13g2_FILL8
XSTDFILL67_1152 VDD VSS sg13g2_FILL8
XSTDFILL67_1160 VDD VSS sg13g2_FILL8
XSTDFILL67_1168 VDD VSS sg13g2_FILL8
XSTDFILL67_1176 VDD VSS sg13g2_FILL8
XSTDFILL67_1184 VDD VSS sg13g2_FILL8
XSTDFILL67_1192 VDD VSS sg13g2_FILL8
XSTDFILL67_1200 VDD VSS sg13g2_FILL8
XSTDFILL67_1208 VDD VSS sg13g2_FILL8
XSTDFILL67_1216 VDD VSS sg13g2_FILL8
XSTDFILL67_1224 VDD VSS sg13g2_FILL8
XSTDFILL67_1232 VDD VSS sg13g2_FILL8
XSTDFILL67_1240 VDD VSS sg13g2_FILL8
XSTDFILL67_1248 VDD VSS sg13g2_FILL8
XSTDFILL67_1256 VDD VSS sg13g2_FILL8
XSTDFILL67_1264 VDD VSS sg13g2_FILL8
XSTDFILL67_1272 VDD VSS sg13g2_FILL8
XSTDFILL67_1280 VDD VSS sg13g2_FILL8
XSTDFILL67_1288 VDD VSS sg13g2_FILL8
XSTDFILL67_1296 VDD VSS sg13g2_FILL8
XSTDFILL67_1304 VDD VSS sg13g2_FILL8
XSTDFILL67_1312 VDD VSS sg13g2_FILL8
XSTDFILL67_1320 VDD VSS sg13g2_FILL8
XSTDFILL67_1328 VDD VSS sg13g2_FILL8
XSTDFILL67_1336 VDD VSS sg13g2_FILL8
XSTDFILL67_1344 VDD VSS sg13g2_FILL8
XSTDFILL67_1352 VDD VSS sg13g2_FILL8
XSTDFILL67_1360 VDD VSS sg13g2_FILL8
XSTDFILL67_1368 VDD VSS sg13g2_FILL8
XSTDFILL67_1376 VDD VSS sg13g2_FILL8
XSTDFILL67_1384 VDD VSS sg13g2_FILL8
XSTDFILL67_1392 VDD VSS sg13g2_FILL8
XSTDFILL67_1400 VDD VSS sg13g2_FILL8
XSTDFILL67_1408 VDD VSS sg13g2_FILL8
XSTDFILL67_1416 VDD VSS sg13g2_FILL8
XSTDFILL67_1424 VDD VSS sg13g2_FILL8
XSTDFILL67_1432 VDD VSS sg13g2_FILL8
XSTDFILL67_1440 VDD VSS sg13g2_FILL8
XSTDFILL67_1448 VDD VSS sg13g2_FILL8
XSTDFILL67_1456 VDD VSS sg13g2_FILL8
XSTDFILL67_1464 VDD VSS sg13g2_FILL8
XSTDFILL67_1472 VDD VSS sg13g2_FILL8
XSTDFILL67_1480 VDD VSS sg13g2_FILL8
XSTDFILL67_1488 VDD VSS sg13g2_FILL8
XSTDFILL67_1496 VDD VSS sg13g2_FILL8
XSTDFILL67_1504 VDD VSS sg13g2_FILL8
XSTDFILL67_1512 VDD VSS sg13g2_FILL8
XSTDFILL67_1520 VDD VSS sg13g2_FILL8
XSTDFILL67_1528 VDD VSS sg13g2_FILL8
XSTDFILL67_1536 VDD VSS sg13g2_FILL8
XSTDFILL67_1544 VDD VSS sg13g2_FILL8
XSTDFILL67_1552 VDD VSS sg13g2_FILL8
XSTDFILL67_1560 VDD VSS sg13g2_FILL8
XSTDFILL67_1568 VDD VSS sg13g2_FILL8
XSTDFILL67_1576 VDD VSS sg13g2_FILL8
XSTDFILL67_1584 VDD VSS sg13g2_FILL8
XSTDFILL67_1592 VDD VSS sg13g2_FILL8
XSTDFILL67_1600 VDD VSS sg13g2_FILL8
XSTDFILL67_1608 VDD VSS sg13g2_FILL8
XSTDFILL67_1616 VDD VSS sg13g2_FILL8
XSTDFILL67_1624 VDD VSS sg13g2_FILL8
XSTDFILL67_1632 VDD VSS sg13g2_FILL8
XSTDFILL67_1640 VDD VSS sg13g2_FILL8
XSTDFILL67_1648 VDD VSS sg13g2_FILL8
XSTDFILL67_1656 VDD VSS sg13g2_FILL8
XSTDFILL67_1664 VDD VSS sg13g2_FILL8
XSTDFILL67_1672 VDD VSS sg13g2_FILL8
XSTDFILL67_1680 VDD VSS sg13g2_FILL8
XSTDFILL67_1688 VDD VSS sg13g2_FILL8
XSTDFILL67_1696 VDD VSS sg13g2_FILL8
XSTDFILL67_1704 VDD VSS sg13g2_FILL8
XSTDFILL67_1712 VDD VSS sg13g2_FILL8
XSTDFILL67_1720 VDD VSS sg13g2_FILL8
XSTDFILL67_1728 VDD VSS sg13g2_FILL8
XSTDFILL67_1736 VDD VSS sg13g2_FILL8
XSTDFILL67_1744 VDD VSS sg13g2_FILL8
XSTDFILL67_1752 VDD VSS sg13g2_FILL8
XSTDFILL67_1760 VDD VSS sg13g2_FILL8
XSTDFILL67_1768 VDD VSS sg13g2_FILL8
XSTDFILL67_1776 VDD VSS sg13g2_FILL8
XSTDFILL67_1784 VDD VSS sg13g2_FILL8
XSTDFILL67_1792 VDD VSS sg13g2_FILL8
XSTDFILL67_1800 VDD VSS sg13g2_FILL8
XSTDFILL67_1808 VDD VSS sg13g2_FILL8
XSTDFILL67_1816 VDD VSS sg13g2_FILL8
XSTDFILL67_1824 VDD VSS sg13g2_FILL8
XSTDFILL67_1832 VDD VSS sg13g2_FILL8
XSTDFILL67_1840 VDD VSS sg13g2_FILL8
XSTDFILL67_1848 VDD VSS sg13g2_FILL8
XSTDFILL67_1856 VDD VSS sg13g2_FILL8
XSTDFILL67_1864 VDD VSS sg13g2_FILL8
XSTDFILL67_1872 VDD VSS sg13g2_FILL8
XSTDFILL67_1880 VDD VSS sg13g2_FILL8
XSTDFILL67_1888 VDD VSS sg13g2_FILL8
XSTDFILL67_1896 VDD VSS sg13g2_FILL8
XSTDFILL67_1904 VDD VSS sg13g2_FILL8
XSTDFILL67_1912 VDD VSS sg13g2_FILL8
XSTDFILL67_1920 VDD VSS sg13g2_FILL8
XSTDFILL67_1928 VDD VSS sg13g2_FILL8
XSTDFILL67_1936 VDD VSS sg13g2_FILL8
XSTDFILL67_1944 VDD VSS sg13g2_FILL8
XSTDFILL67_1952 VDD VSS sg13g2_FILL8
XSTDFILL67_1960 VDD VSS sg13g2_FILL8
XSTDFILL67_1968 VDD VSS sg13g2_FILL8
XSTDFILL67_1976 VDD VSS sg13g2_FILL8
XSTDFILL67_1984 VDD VSS sg13g2_FILL8
XSTDFILL67_1992 VDD VSS sg13g2_FILL8
XSTDFILL67_2000 VDD VSS sg13g2_FILL8
XSTDFILL67_2008 VDD VSS sg13g2_FILL8
XSTDFILL67_2016 VDD VSS sg13g2_FILL8
XSTDFILL67_2024 VDD VSS sg13g2_FILL8
XSTDFILL67_2032 VDD VSS sg13g2_FILL8
XSTDFILL67_2040 VDD VSS sg13g2_FILL8
XSTDFILL67_2048 VDD VSS sg13g2_FILL8
XSTDFILL67_2056 VDD VSS sg13g2_FILL8
XSTDFILL67_2064 VDD VSS sg13g2_FILL8
XSTDFILL67_2072 VDD VSS sg13g2_FILL8
XSTDFILL67_2080 VDD VSS sg13g2_FILL8
XSTDFILL67_2088 VDD VSS sg13g2_FILL8
XSTDFILL67_2096 VDD VSS sg13g2_FILL8
XSTDFILL67_2104 VDD VSS sg13g2_FILL8
XSTDFILL67_2112 VDD VSS sg13g2_FILL8
XSTDFILL67_2120 VDD VSS sg13g2_FILL8
XSTDFILL67_2128 VDD VSS sg13g2_FILL8
XSTDFILL67_2136 VDD VSS sg13g2_FILL8
XSTDFILL67_2144 VDD VSS sg13g2_FILL8
XSTDFILL67_2152 VDD VSS sg13g2_FILL8
XSTDFILL67_2160 VDD VSS sg13g2_FILL8
XSTDFILL67_2168 VDD VSS sg13g2_FILL4
XSTDFILL68_0 VDD VSS sg13g2_FILL8
XSTDFILL68_8 VDD VSS sg13g2_FILL8
XSTDFILL68_16 VDD VSS sg13g2_FILL8
XSTDFILL68_24 VDD VSS sg13g2_FILL8
XSTDFILL68_32 VDD VSS sg13g2_FILL8
XSTDFILL68_40 VDD VSS sg13g2_FILL8
XSTDFILL68_48 VDD VSS sg13g2_FILL8
XSTDFILL68_56 VDD VSS sg13g2_FILL8
XSTDFILL68_64 VDD VSS sg13g2_FILL8
XSTDFILL68_72 VDD VSS sg13g2_FILL8
XSTDFILL68_80 VDD VSS sg13g2_FILL8
XSTDFILL68_88 VDD VSS sg13g2_FILL8
XSTDFILL68_96 VDD VSS sg13g2_FILL8
XSTDFILL68_104 VDD VSS sg13g2_FILL8
XSTDFILL68_112 VDD VSS sg13g2_FILL8
XSTDFILL68_120 VDD VSS sg13g2_FILL8
XSTDFILL68_128 VDD VSS sg13g2_FILL8
XSTDFILL68_136 VDD VSS sg13g2_FILL8
XSTDFILL68_144 VDD VSS sg13g2_FILL8
XSTDFILL68_152 VDD VSS sg13g2_FILL8
XSTDFILL68_160 VDD VSS sg13g2_FILL8
XSTDFILL68_168 VDD VSS sg13g2_FILL8
XSTDFILL68_176 VDD VSS sg13g2_FILL8
XSTDFILL68_184 VDD VSS sg13g2_FILL8
XSTDFILL68_192 VDD VSS sg13g2_FILL8
XSTDFILL68_200 VDD VSS sg13g2_FILL8
XSTDFILL68_208 VDD VSS sg13g2_FILL8
XSTDFILL68_216 VDD VSS sg13g2_FILL8
XSTDFILL68_224 VDD VSS sg13g2_FILL8
XSTDFILL68_232 VDD VSS sg13g2_FILL8
XSTDFILL68_240 VDD VSS sg13g2_FILL8
XSTDFILL68_248 VDD VSS sg13g2_FILL8
XSTDFILL68_256 VDD VSS sg13g2_FILL8
XSTDFILL68_264 VDD VSS sg13g2_FILL8
XSTDFILL68_272 VDD VSS sg13g2_FILL8
XSTDFILL68_280 VDD VSS sg13g2_FILL8
XSTDFILL68_288 VDD VSS sg13g2_FILL8
XSTDFILL68_296 VDD VSS sg13g2_FILL8
XSTDFILL68_304 VDD VSS sg13g2_FILL8
XSTDFILL68_312 VDD VSS sg13g2_FILL8
XSTDFILL68_320 VDD VSS sg13g2_FILL8
XSTDFILL68_328 VDD VSS sg13g2_FILL8
XSTDFILL68_336 VDD VSS sg13g2_FILL8
XSTDFILL68_344 VDD VSS sg13g2_FILL8
XSTDFILL68_352 VDD VSS sg13g2_FILL8
XSTDFILL68_360 VDD VSS sg13g2_FILL8
XSTDFILL68_368 VDD VSS sg13g2_FILL8
XSTDFILL68_376 VDD VSS sg13g2_FILL8
XSTDFILL68_384 VDD VSS sg13g2_FILL8
XSTDFILL68_392 VDD VSS sg13g2_FILL8
XSTDFILL68_400 VDD VSS sg13g2_FILL8
XSTDFILL68_408 VDD VSS sg13g2_FILL8
XSTDFILL68_416 VDD VSS sg13g2_FILL8
XSTDFILL68_424 VDD VSS sg13g2_FILL8
XSTDFILL68_432 VDD VSS sg13g2_FILL8
XSTDFILL68_440 VDD VSS sg13g2_FILL8
XSTDFILL68_448 VDD VSS sg13g2_FILL8
XSTDFILL68_456 VDD VSS sg13g2_FILL8
XSTDFILL68_464 VDD VSS sg13g2_FILL8
XSTDFILL68_472 VDD VSS sg13g2_FILL8
XSTDFILL68_480 VDD VSS sg13g2_FILL8
XSTDFILL68_488 VDD VSS sg13g2_FILL8
XSTDFILL68_496 VDD VSS sg13g2_FILL8
XSTDFILL68_504 VDD VSS sg13g2_FILL8
XSTDFILL68_512 VDD VSS sg13g2_FILL8
XSTDFILL68_520 VDD VSS sg13g2_FILL8
XSTDFILL68_528 VDD VSS sg13g2_FILL8
XSTDFILL68_536 VDD VSS sg13g2_FILL8
XSTDFILL68_544 VDD VSS sg13g2_FILL8
XSTDFILL68_552 VDD VSS sg13g2_FILL8
XSTDFILL68_560 VDD VSS sg13g2_FILL8
XSTDFILL68_568 VDD VSS sg13g2_FILL8
XSTDFILL68_576 VDD VSS sg13g2_FILL8
XSTDFILL68_584 VDD VSS sg13g2_FILL8
XSTDFILL68_592 VDD VSS sg13g2_FILL8
XSTDFILL68_600 VDD VSS sg13g2_FILL8
XSTDFILL68_608 VDD VSS sg13g2_FILL8
XSTDFILL68_616 VDD VSS sg13g2_FILL8
XSTDFILL68_624 VDD VSS sg13g2_FILL8
XSTDFILL68_632 VDD VSS sg13g2_FILL8
XSTDFILL68_640 VDD VSS sg13g2_FILL8
XSTDFILL68_648 VDD VSS sg13g2_FILL8
XSTDFILL68_656 VDD VSS sg13g2_FILL8
XSTDFILL68_664 VDD VSS sg13g2_FILL8
XSTDFILL68_672 VDD VSS sg13g2_FILL8
XSTDFILL68_680 VDD VSS sg13g2_FILL8
XSTDFILL68_688 VDD VSS sg13g2_FILL8
XSTDFILL68_696 VDD VSS sg13g2_FILL8
XSTDFILL68_704 VDD VSS sg13g2_FILL8
XSTDFILL68_712 VDD VSS sg13g2_FILL8
XSTDFILL68_720 VDD VSS sg13g2_FILL8
XSTDFILL68_728 VDD VSS sg13g2_FILL8
XSTDFILL68_736 VDD VSS sg13g2_FILL8
XSTDFILL68_744 VDD VSS sg13g2_FILL8
XSTDFILL68_752 VDD VSS sg13g2_FILL8
XSTDFILL68_760 VDD VSS sg13g2_FILL8
XSTDFILL68_768 VDD VSS sg13g2_FILL8
XSTDFILL68_776 VDD VSS sg13g2_FILL8
XSTDFILL68_784 VDD VSS sg13g2_FILL8
XSTDFILL68_792 VDD VSS sg13g2_FILL8
XSTDFILL68_800 VDD VSS sg13g2_FILL8
XSTDFILL68_808 VDD VSS sg13g2_FILL8
XSTDFILL68_816 VDD VSS sg13g2_FILL8
XSTDFILL68_824 VDD VSS sg13g2_FILL8
XSTDFILL68_832 VDD VSS sg13g2_FILL8
XSTDFILL68_840 VDD VSS sg13g2_FILL8
XSTDFILL68_848 VDD VSS sg13g2_FILL8
XSTDFILL68_856 VDD VSS sg13g2_FILL8
XSTDFILL68_864 VDD VSS sg13g2_FILL8
XSTDFILL68_872 VDD VSS sg13g2_FILL8
XSTDFILL68_880 VDD VSS sg13g2_FILL8
XSTDFILL68_888 VDD VSS sg13g2_FILL8
XSTDFILL68_896 VDD VSS sg13g2_FILL8
XSTDFILL68_904 VDD VSS sg13g2_FILL8
XSTDFILL68_912 VDD VSS sg13g2_FILL8
XSTDFILL68_920 VDD VSS sg13g2_FILL8
XSTDFILL68_928 VDD VSS sg13g2_FILL8
XSTDFILL68_936 VDD VSS sg13g2_FILL8
XSTDFILL68_944 VDD VSS sg13g2_FILL8
XSTDFILL68_952 VDD VSS sg13g2_FILL8
XSTDFILL68_960 VDD VSS sg13g2_FILL8
XSTDFILL68_968 VDD VSS sg13g2_FILL8
XSTDFILL68_976 VDD VSS sg13g2_FILL8
XSTDFILL68_984 VDD VSS sg13g2_FILL8
XSTDFILL68_992 VDD VSS sg13g2_FILL8
XSTDFILL68_1000 VDD VSS sg13g2_FILL8
XSTDFILL68_1008 VDD VSS sg13g2_FILL8
XSTDFILL68_1016 VDD VSS sg13g2_FILL8
XSTDFILL68_1024 VDD VSS sg13g2_FILL8
XSTDFILL68_1032 VDD VSS sg13g2_FILL8
XSTDFILL68_1040 VDD VSS sg13g2_FILL8
XSTDFILL68_1048 VDD VSS sg13g2_FILL8
XSTDFILL68_1056 VDD VSS sg13g2_FILL8
XSTDFILL68_1064 VDD VSS sg13g2_FILL8
XSTDFILL68_1072 VDD VSS sg13g2_FILL8
XSTDFILL68_1080 VDD VSS sg13g2_FILL8
XSTDFILL68_1088 VDD VSS sg13g2_FILL8
XSTDFILL68_1096 VDD VSS sg13g2_FILL8
XSTDFILL68_1104 VDD VSS sg13g2_FILL8
XSTDFILL68_1112 VDD VSS sg13g2_FILL8
XSTDFILL68_1120 VDD VSS sg13g2_FILL8
XSTDFILL68_1128 VDD VSS sg13g2_FILL8
XSTDFILL68_1136 VDD VSS sg13g2_FILL8
XSTDFILL68_1144 VDD VSS sg13g2_FILL8
XSTDFILL68_1152 VDD VSS sg13g2_FILL8
XSTDFILL68_1160 VDD VSS sg13g2_FILL8
XSTDFILL68_1168 VDD VSS sg13g2_FILL8
XSTDFILL68_1176 VDD VSS sg13g2_FILL8
XSTDFILL68_1184 VDD VSS sg13g2_FILL8
XSTDFILL68_1192 VDD VSS sg13g2_FILL8
XSTDFILL68_1200 VDD VSS sg13g2_FILL8
XSTDFILL68_1208 VDD VSS sg13g2_FILL8
XSTDFILL68_1216 VDD VSS sg13g2_FILL8
XSTDFILL68_1224 VDD VSS sg13g2_FILL8
XSTDFILL68_1232 VDD VSS sg13g2_FILL8
XSTDFILL68_1240 VDD VSS sg13g2_FILL8
XSTDFILL68_1248 VDD VSS sg13g2_FILL8
XSTDFILL68_1256 VDD VSS sg13g2_FILL8
XSTDFILL68_1264 VDD VSS sg13g2_FILL8
XSTDFILL68_1272 VDD VSS sg13g2_FILL8
XSTDFILL68_1280 VDD VSS sg13g2_FILL8
XSTDFILL68_1288 VDD VSS sg13g2_FILL8
XSTDFILL68_1296 VDD VSS sg13g2_FILL8
XSTDFILL68_1304 VDD VSS sg13g2_FILL8
XSTDFILL68_1312 VDD VSS sg13g2_FILL8
XSTDFILL68_1320 VDD VSS sg13g2_FILL8
XSTDFILL68_1328 VDD VSS sg13g2_FILL8
XSTDFILL68_1336 VDD VSS sg13g2_FILL8
XSTDFILL68_1344 VDD VSS sg13g2_FILL8
XSTDFILL68_1352 VDD VSS sg13g2_FILL8
XSTDFILL68_1360 VDD VSS sg13g2_FILL8
XSTDFILL68_1368 VDD VSS sg13g2_FILL8
XSTDFILL68_1376 VDD VSS sg13g2_FILL8
XSTDFILL68_1384 VDD VSS sg13g2_FILL8
XSTDFILL68_1392 VDD VSS sg13g2_FILL8
XSTDFILL68_1400 VDD VSS sg13g2_FILL8
XSTDFILL68_1408 VDD VSS sg13g2_FILL8
XSTDFILL68_1416 VDD VSS sg13g2_FILL8
XSTDFILL68_1424 VDD VSS sg13g2_FILL8
XSTDFILL68_1432 VDD VSS sg13g2_FILL8
XSTDFILL68_1440 VDD VSS sg13g2_FILL8
XSTDFILL68_1448 VDD VSS sg13g2_FILL8
XSTDFILL68_1456 VDD VSS sg13g2_FILL8
XSTDFILL68_1464 VDD VSS sg13g2_FILL8
XSTDFILL68_1472 VDD VSS sg13g2_FILL8
XSTDFILL68_1480 VDD VSS sg13g2_FILL8
XSTDFILL68_1488 VDD VSS sg13g2_FILL8
XSTDFILL68_1496 VDD VSS sg13g2_FILL8
XSTDFILL68_1504 VDD VSS sg13g2_FILL8
XSTDFILL68_1512 VDD VSS sg13g2_FILL8
XSTDFILL68_1520 VDD VSS sg13g2_FILL8
XSTDFILL68_1528 VDD VSS sg13g2_FILL8
XSTDFILL68_1536 VDD VSS sg13g2_FILL8
XSTDFILL68_1544 VDD VSS sg13g2_FILL8
XSTDFILL68_1552 VDD VSS sg13g2_FILL8
XSTDFILL68_1560 VDD VSS sg13g2_FILL8
XSTDFILL68_1568 VDD VSS sg13g2_FILL8
XSTDFILL68_1576 VDD VSS sg13g2_FILL8
XSTDFILL68_1584 VDD VSS sg13g2_FILL8
XSTDFILL68_1592 VDD VSS sg13g2_FILL8
XSTDFILL68_1600 VDD VSS sg13g2_FILL8
XSTDFILL68_1608 VDD VSS sg13g2_FILL8
XSTDFILL68_1616 VDD VSS sg13g2_FILL8
XSTDFILL68_1624 VDD VSS sg13g2_FILL8
XSTDFILL68_1632 VDD VSS sg13g2_FILL8
XSTDFILL68_1640 VDD VSS sg13g2_FILL8
XSTDFILL68_1648 VDD VSS sg13g2_FILL8
XSTDFILL68_1656 VDD VSS sg13g2_FILL8
XSTDFILL68_1664 VDD VSS sg13g2_FILL8
XSTDFILL68_1672 VDD VSS sg13g2_FILL8
XSTDFILL68_1680 VDD VSS sg13g2_FILL8
XSTDFILL68_1688 VDD VSS sg13g2_FILL8
XSTDFILL68_1696 VDD VSS sg13g2_FILL8
XSTDFILL68_1704 VDD VSS sg13g2_FILL8
XSTDFILL68_1712 VDD VSS sg13g2_FILL8
XSTDFILL68_1720 VDD VSS sg13g2_FILL8
XSTDFILL68_1728 VDD VSS sg13g2_FILL8
XSTDFILL68_1736 VDD VSS sg13g2_FILL8
XSTDFILL68_1744 VDD VSS sg13g2_FILL8
XSTDFILL68_1752 VDD VSS sg13g2_FILL8
XSTDFILL68_1760 VDD VSS sg13g2_FILL8
XSTDFILL68_1768 VDD VSS sg13g2_FILL8
XSTDFILL68_1776 VDD VSS sg13g2_FILL8
XSTDFILL68_1784 VDD VSS sg13g2_FILL8
XSTDFILL68_1792 VDD VSS sg13g2_FILL8
XSTDFILL68_1800 VDD VSS sg13g2_FILL8
XSTDFILL68_1808 VDD VSS sg13g2_FILL8
XSTDFILL68_1816 VDD VSS sg13g2_FILL8
XSTDFILL68_1824 VDD VSS sg13g2_FILL8
XSTDFILL68_1832 VDD VSS sg13g2_FILL8
XSTDFILL68_1840 VDD VSS sg13g2_FILL8
XSTDFILL68_1848 VDD VSS sg13g2_FILL8
XSTDFILL68_1856 VDD VSS sg13g2_FILL8
XSTDFILL68_1864 VDD VSS sg13g2_FILL8
XSTDFILL68_1872 VDD VSS sg13g2_FILL8
XSTDFILL68_1880 VDD VSS sg13g2_FILL8
XSTDFILL68_1888 VDD VSS sg13g2_FILL8
XSTDFILL68_1896 VDD VSS sg13g2_FILL8
XSTDFILL68_1904 VDD VSS sg13g2_FILL8
XSTDFILL68_1912 VDD VSS sg13g2_FILL8
XSTDFILL68_1920 VDD VSS sg13g2_FILL8
XSTDFILL68_1928 VDD VSS sg13g2_FILL8
XSTDFILL68_1936 VDD VSS sg13g2_FILL8
XSTDFILL68_1944 VDD VSS sg13g2_FILL8
XSTDFILL68_1952 VDD VSS sg13g2_FILL8
XSTDFILL68_1960 VDD VSS sg13g2_FILL8
XSTDFILL68_1968 VDD VSS sg13g2_FILL8
XSTDFILL68_1976 VDD VSS sg13g2_FILL8
XSTDFILL68_1984 VDD VSS sg13g2_FILL8
XSTDFILL68_1992 VDD VSS sg13g2_FILL8
XSTDFILL68_2000 VDD VSS sg13g2_FILL8
XSTDFILL68_2008 VDD VSS sg13g2_FILL8
XSTDFILL68_2016 VDD VSS sg13g2_FILL8
XSTDFILL68_2024 VDD VSS sg13g2_FILL8
XSTDFILL68_2032 VDD VSS sg13g2_FILL8
XSTDFILL68_2040 VDD VSS sg13g2_FILL8
XSTDFILL68_2048 VDD VSS sg13g2_FILL8
XSTDFILL68_2056 VDD VSS sg13g2_FILL8
XSTDFILL68_2064 VDD VSS sg13g2_FILL8
XSTDFILL68_2072 VDD VSS sg13g2_FILL8
XSTDFILL68_2080 VDD VSS sg13g2_FILL8
XSTDFILL68_2088 VDD VSS sg13g2_FILL8
XSTDFILL68_2096 VDD VSS sg13g2_FILL8
XSTDFILL68_2104 VDD VSS sg13g2_FILL8
XSTDFILL68_2112 VDD VSS sg13g2_FILL8
XSTDFILL68_2120 VDD VSS sg13g2_FILL8
XSTDFILL68_2128 VDD VSS sg13g2_FILL8
XSTDFILL68_2136 VDD VSS sg13g2_FILL8
XSTDFILL68_2144 VDD VSS sg13g2_FILL8
XSTDFILL68_2152 VDD VSS sg13g2_FILL8
XSTDFILL68_2160 VDD VSS sg13g2_FILL8
XSTDFILL68_2168 VDD VSS sg13g2_FILL4
XSTDFILL69_0 VDD VSS sg13g2_FILL8
XSTDFILL69_8 VDD VSS sg13g2_FILL8
XSTDFILL69_16 VDD VSS sg13g2_FILL8
XSTDFILL69_24 VDD VSS sg13g2_FILL8
XSTDFILL69_32 VDD VSS sg13g2_FILL8
XSTDFILL69_40 VDD VSS sg13g2_FILL8
XSTDFILL69_48 VDD VSS sg13g2_FILL8
XSTDFILL69_56 VDD VSS sg13g2_FILL8
XSTDFILL69_64 VDD VSS sg13g2_FILL8
XSTDFILL69_72 VDD VSS sg13g2_FILL8
XSTDFILL69_80 VDD VSS sg13g2_FILL8
XSTDFILL69_88 VDD VSS sg13g2_FILL8
XSTDFILL69_96 VDD VSS sg13g2_FILL8
XSTDFILL69_104 VDD VSS sg13g2_FILL8
XSTDFILL69_112 VDD VSS sg13g2_FILL8
XSTDFILL69_120 VDD VSS sg13g2_FILL8
XSTDFILL69_128 VDD VSS sg13g2_FILL8
XSTDFILL69_136 VDD VSS sg13g2_FILL8
XSTDFILL69_144 VDD VSS sg13g2_FILL8
XSTDFILL69_152 VDD VSS sg13g2_FILL8
XSTDFILL69_160 VDD VSS sg13g2_FILL8
XSTDFILL69_168 VDD VSS sg13g2_FILL8
XSTDFILL69_176 VDD VSS sg13g2_FILL8
XSTDFILL69_184 VDD VSS sg13g2_FILL8
XSTDFILL69_192 VDD VSS sg13g2_FILL8
XSTDFILL69_200 VDD VSS sg13g2_FILL8
XSTDFILL69_208 VDD VSS sg13g2_FILL8
XSTDFILL69_216 VDD VSS sg13g2_FILL8
XSTDFILL69_224 VDD VSS sg13g2_FILL8
XSTDFILL69_232 VDD VSS sg13g2_FILL8
XSTDFILL69_240 VDD VSS sg13g2_FILL8
XSTDFILL69_248 VDD VSS sg13g2_FILL8
XSTDFILL69_256 VDD VSS sg13g2_FILL8
XSTDFILL69_264 VDD VSS sg13g2_FILL8
XSTDFILL69_272 VDD VSS sg13g2_FILL8
XSTDFILL69_280 VDD VSS sg13g2_FILL8
XSTDFILL69_288 VDD VSS sg13g2_FILL8
XSTDFILL69_296 VDD VSS sg13g2_FILL8
XSTDFILL69_304 VDD VSS sg13g2_FILL8
XSTDFILL69_312 VDD VSS sg13g2_FILL8
XSTDFILL69_320 VDD VSS sg13g2_FILL8
XSTDFILL69_328 VDD VSS sg13g2_FILL8
XSTDFILL69_336 VDD VSS sg13g2_FILL8
XSTDFILL69_344 VDD VSS sg13g2_FILL8
XSTDFILL69_352 VDD VSS sg13g2_FILL8
XSTDFILL69_360 VDD VSS sg13g2_FILL8
XSTDFILL69_368 VDD VSS sg13g2_FILL8
XSTDFILL69_376 VDD VSS sg13g2_FILL8
XSTDFILL69_384 VDD VSS sg13g2_FILL8
XSTDFILL69_392 VDD VSS sg13g2_FILL8
XSTDFILL69_400 VDD VSS sg13g2_FILL8
XSTDFILL69_408 VDD VSS sg13g2_FILL8
XSTDFILL69_416 VDD VSS sg13g2_FILL8
XSTDFILL69_424 VDD VSS sg13g2_FILL8
XSTDFILL69_432 VDD VSS sg13g2_FILL8
XSTDFILL69_440 VDD VSS sg13g2_FILL8
XSTDFILL69_448 VDD VSS sg13g2_FILL8
XSTDFILL69_456 VDD VSS sg13g2_FILL8
XSTDFILL69_464 VDD VSS sg13g2_FILL8
XSTDFILL69_472 VDD VSS sg13g2_FILL8
XSTDFILL69_480 VDD VSS sg13g2_FILL8
XSTDFILL69_488 VDD VSS sg13g2_FILL8
XSTDFILL69_496 VDD VSS sg13g2_FILL8
XSTDFILL69_504 VDD VSS sg13g2_FILL8
XSTDFILL69_512 VDD VSS sg13g2_FILL8
XSTDFILL69_520 VDD VSS sg13g2_FILL8
XSTDFILL69_528 VDD VSS sg13g2_FILL8
XSTDFILL69_536 VDD VSS sg13g2_FILL8
XSTDFILL69_544 VDD VSS sg13g2_FILL8
XSTDFILL69_552 VDD VSS sg13g2_FILL8
XSTDFILL69_560 VDD VSS sg13g2_FILL8
XSTDFILL69_568 VDD VSS sg13g2_FILL8
XSTDFILL69_576 VDD VSS sg13g2_FILL8
XSTDFILL69_584 VDD VSS sg13g2_FILL8
XSTDFILL69_592 VDD VSS sg13g2_FILL8
XSTDFILL69_600 VDD VSS sg13g2_FILL8
XSTDFILL69_608 VDD VSS sg13g2_FILL8
XSTDFILL69_616 VDD VSS sg13g2_FILL8
XSTDFILL69_624 VDD VSS sg13g2_FILL8
XSTDFILL69_632 VDD VSS sg13g2_FILL8
XSTDFILL69_640 VDD VSS sg13g2_FILL8
XSTDFILL69_648 VDD VSS sg13g2_FILL8
XSTDFILL69_656 VDD VSS sg13g2_FILL8
XSTDFILL69_664 VDD VSS sg13g2_FILL8
XSTDFILL69_672 VDD VSS sg13g2_FILL8
XSTDFILL69_680 VDD VSS sg13g2_FILL8
XSTDFILL69_688 VDD VSS sg13g2_FILL8
XSTDFILL69_696 VDD VSS sg13g2_FILL8
XSTDFILL69_704 VDD VSS sg13g2_FILL8
XSTDFILL69_712 VDD VSS sg13g2_FILL8
XSTDFILL69_720 VDD VSS sg13g2_FILL8
XSTDFILL69_728 VDD VSS sg13g2_FILL8
XSTDFILL69_736 VDD VSS sg13g2_FILL8
XSTDFILL69_744 VDD VSS sg13g2_FILL8
XSTDFILL69_752 VDD VSS sg13g2_FILL8
XSTDFILL69_760 VDD VSS sg13g2_FILL8
XSTDFILL69_768 VDD VSS sg13g2_FILL8
XSTDFILL69_776 VDD VSS sg13g2_FILL8
XSTDFILL69_784 VDD VSS sg13g2_FILL8
XSTDFILL69_792 VDD VSS sg13g2_FILL8
XSTDFILL69_800 VDD VSS sg13g2_FILL8
XSTDFILL69_808 VDD VSS sg13g2_FILL8
XSTDFILL69_816 VDD VSS sg13g2_FILL8
XSTDFILL69_824 VDD VSS sg13g2_FILL8
XSTDFILL69_832 VDD VSS sg13g2_FILL8
XSTDFILL69_840 VDD VSS sg13g2_FILL8
XSTDFILL69_848 VDD VSS sg13g2_FILL8
XSTDFILL69_856 VDD VSS sg13g2_FILL8
XSTDFILL69_864 VDD VSS sg13g2_FILL8
XSTDFILL69_872 VDD VSS sg13g2_FILL8
XSTDFILL69_880 VDD VSS sg13g2_FILL8
XSTDFILL69_888 VDD VSS sg13g2_FILL8
XSTDFILL69_896 VDD VSS sg13g2_FILL8
XSTDFILL69_904 VDD VSS sg13g2_FILL8
XSTDFILL69_912 VDD VSS sg13g2_FILL8
XSTDFILL69_920 VDD VSS sg13g2_FILL8
XSTDFILL69_928 VDD VSS sg13g2_FILL8
XSTDFILL69_936 VDD VSS sg13g2_FILL8
XSTDFILL69_944 VDD VSS sg13g2_FILL8
XSTDFILL69_952 VDD VSS sg13g2_FILL8
XSTDFILL69_960 VDD VSS sg13g2_FILL8
XSTDFILL69_968 VDD VSS sg13g2_FILL8
XSTDFILL69_976 VDD VSS sg13g2_FILL8
XSTDFILL69_984 VDD VSS sg13g2_FILL8
XSTDFILL69_992 VDD VSS sg13g2_FILL8
XSTDFILL69_1000 VDD VSS sg13g2_FILL8
XSTDFILL69_1008 VDD VSS sg13g2_FILL8
XSTDFILL69_1016 VDD VSS sg13g2_FILL8
XSTDFILL69_1024 VDD VSS sg13g2_FILL8
XSTDFILL69_1032 VDD VSS sg13g2_FILL8
XSTDFILL69_1040 VDD VSS sg13g2_FILL8
XSTDFILL69_1048 VDD VSS sg13g2_FILL8
XSTDFILL69_1056 VDD VSS sg13g2_FILL8
XSTDFILL69_1064 VDD VSS sg13g2_FILL8
XSTDFILL69_1072 VDD VSS sg13g2_FILL8
XSTDFILL69_1080 VDD VSS sg13g2_FILL8
XSTDFILL69_1088 VDD VSS sg13g2_FILL8
XSTDFILL69_1096 VDD VSS sg13g2_FILL8
XSTDFILL69_1104 VDD VSS sg13g2_FILL8
XSTDFILL69_1112 VDD VSS sg13g2_FILL8
XSTDFILL69_1120 VDD VSS sg13g2_FILL8
XSTDFILL69_1128 VDD VSS sg13g2_FILL8
XSTDFILL69_1136 VDD VSS sg13g2_FILL8
XSTDFILL69_1144 VDD VSS sg13g2_FILL8
XSTDFILL69_1152 VDD VSS sg13g2_FILL8
XSTDFILL69_1160 VDD VSS sg13g2_FILL8
XSTDFILL69_1168 VDD VSS sg13g2_FILL8
XSTDFILL69_1176 VDD VSS sg13g2_FILL8
XSTDFILL69_1184 VDD VSS sg13g2_FILL8
XSTDFILL69_1192 VDD VSS sg13g2_FILL8
XSTDFILL69_1200 VDD VSS sg13g2_FILL8
XSTDFILL69_1208 VDD VSS sg13g2_FILL8
XSTDFILL69_1216 VDD VSS sg13g2_FILL8
XSTDFILL69_1224 VDD VSS sg13g2_FILL8
XSTDFILL69_1232 VDD VSS sg13g2_FILL8
XSTDFILL69_1240 VDD VSS sg13g2_FILL8
XSTDFILL69_1248 VDD VSS sg13g2_FILL8
XSTDFILL69_1256 VDD VSS sg13g2_FILL8
XSTDFILL69_1264 VDD VSS sg13g2_FILL8
XSTDFILL69_1272 VDD VSS sg13g2_FILL8
XSTDFILL69_1280 VDD VSS sg13g2_FILL8
XSTDFILL69_1288 VDD VSS sg13g2_FILL8
XSTDFILL69_1296 VDD VSS sg13g2_FILL8
XSTDFILL69_1304 VDD VSS sg13g2_FILL8
XSTDFILL69_1312 VDD VSS sg13g2_FILL8
XSTDFILL69_1320 VDD VSS sg13g2_FILL8
XSTDFILL69_1328 VDD VSS sg13g2_FILL8
XSTDFILL69_1336 VDD VSS sg13g2_FILL8
XSTDFILL69_1344 VDD VSS sg13g2_FILL8
XSTDFILL69_1352 VDD VSS sg13g2_FILL8
XSTDFILL69_1360 VDD VSS sg13g2_FILL8
XSTDFILL69_1368 VDD VSS sg13g2_FILL8
XSTDFILL69_1376 VDD VSS sg13g2_FILL8
XSTDFILL69_1384 VDD VSS sg13g2_FILL8
XSTDFILL69_1392 VDD VSS sg13g2_FILL8
XSTDFILL69_1400 VDD VSS sg13g2_FILL8
XSTDFILL69_1408 VDD VSS sg13g2_FILL8
XSTDFILL69_1416 VDD VSS sg13g2_FILL8
XSTDFILL69_1424 VDD VSS sg13g2_FILL8
XSTDFILL69_1432 VDD VSS sg13g2_FILL8
XSTDFILL69_1440 VDD VSS sg13g2_FILL8
XSTDFILL69_1448 VDD VSS sg13g2_FILL8
XSTDFILL69_1456 VDD VSS sg13g2_FILL8
XSTDFILL69_1464 VDD VSS sg13g2_FILL8
XSTDFILL69_1472 VDD VSS sg13g2_FILL8
XSTDFILL69_1480 VDD VSS sg13g2_FILL8
XSTDFILL69_1488 VDD VSS sg13g2_FILL8
XSTDFILL69_1496 VDD VSS sg13g2_FILL8
XSTDFILL69_1504 VDD VSS sg13g2_FILL8
XSTDFILL69_1512 VDD VSS sg13g2_FILL8
XSTDFILL69_1520 VDD VSS sg13g2_FILL8
XSTDFILL69_1528 VDD VSS sg13g2_FILL8
XSTDFILL69_1536 VDD VSS sg13g2_FILL8
XSTDFILL69_1544 VDD VSS sg13g2_FILL8
XSTDFILL69_1552 VDD VSS sg13g2_FILL8
XSTDFILL69_1560 VDD VSS sg13g2_FILL8
XSTDFILL69_1568 VDD VSS sg13g2_FILL8
XSTDFILL69_1576 VDD VSS sg13g2_FILL8
XSTDFILL69_1584 VDD VSS sg13g2_FILL8
XSTDFILL69_1592 VDD VSS sg13g2_FILL8
XSTDFILL69_1600 VDD VSS sg13g2_FILL8
XSTDFILL69_1608 VDD VSS sg13g2_FILL8
XSTDFILL69_1616 VDD VSS sg13g2_FILL8
XSTDFILL69_1624 VDD VSS sg13g2_FILL8
XSTDFILL69_1632 VDD VSS sg13g2_FILL8
XSTDFILL69_1640 VDD VSS sg13g2_FILL8
XSTDFILL69_1648 VDD VSS sg13g2_FILL8
XSTDFILL69_1656 VDD VSS sg13g2_FILL8
XSTDFILL69_1664 VDD VSS sg13g2_FILL8
XSTDFILL69_1672 VDD VSS sg13g2_FILL8
XSTDFILL69_1680 VDD VSS sg13g2_FILL8
XSTDFILL69_1688 VDD VSS sg13g2_FILL8
XSTDFILL69_1696 VDD VSS sg13g2_FILL8
XSTDFILL69_1704 VDD VSS sg13g2_FILL8
XSTDFILL69_1712 VDD VSS sg13g2_FILL8
XSTDFILL69_1720 VDD VSS sg13g2_FILL8
XSTDFILL69_1728 VDD VSS sg13g2_FILL8
XSTDFILL69_1736 VDD VSS sg13g2_FILL8
XSTDFILL69_1744 VDD VSS sg13g2_FILL8
XSTDFILL69_1752 VDD VSS sg13g2_FILL8
XSTDFILL69_1760 VDD VSS sg13g2_FILL8
XSTDFILL69_1768 VDD VSS sg13g2_FILL8
XSTDFILL69_1776 VDD VSS sg13g2_FILL8
XSTDFILL69_1784 VDD VSS sg13g2_FILL8
XSTDFILL69_1792 VDD VSS sg13g2_FILL8
XSTDFILL69_1800 VDD VSS sg13g2_FILL8
XSTDFILL69_1808 VDD VSS sg13g2_FILL8
XSTDFILL69_1816 VDD VSS sg13g2_FILL8
XSTDFILL69_1824 VDD VSS sg13g2_FILL8
XSTDFILL69_1832 VDD VSS sg13g2_FILL8
XSTDFILL69_1840 VDD VSS sg13g2_FILL8
XSTDFILL69_1848 VDD VSS sg13g2_FILL8
XSTDFILL69_1856 VDD VSS sg13g2_FILL8
XSTDFILL69_1864 VDD VSS sg13g2_FILL8
XSTDFILL69_1872 VDD VSS sg13g2_FILL8
XSTDFILL69_1880 VDD VSS sg13g2_FILL8
XSTDFILL69_1888 VDD VSS sg13g2_FILL8
XSTDFILL69_1896 VDD VSS sg13g2_FILL8
XSTDFILL69_1904 VDD VSS sg13g2_FILL8
XSTDFILL69_1912 VDD VSS sg13g2_FILL8
XSTDFILL69_1920 VDD VSS sg13g2_FILL8
XSTDFILL69_1928 VDD VSS sg13g2_FILL8
XSTDFILL69_1936 VDD VSS sg13g2_FILL8
XSTDFILL69_1944 VDD VSS sg13g2_FILL8
XSTDFILL69_1952 VDD VSS sg13g2_FILL8
XSTDFILL69_1960 VDD VSS sg13g2_FILL8
XSTDFILL69_1968 VDD VSS sg13g2_FILL8
XSTDFILL69_1976 VDD VSS sg13g2_FILL8
XSTDFILL69_1984 VDD VSS sg13g2_FILL8
XSTDFILL69_1992 VDD VSS sg13g2_FILL8
XSTDFILL69_2000 VDD VSS sg13g2_FILL8
XSTDFILL69_2008 VDD VSS sg13g2_FILL8
XSTDFILL69_2016 VDD VSS sg13g2_FILL8
XSTDFILL69_2024 VDD VSS sg13g2_FILL8
XSTDFILL69_2032 VDD VSS sg13g2_FILL8
XSTDFILL69_2040 VDD VSS sg13g2_FILL8
XSTDFILL69_2048 VDD VSS sg13g2_FILL8
XSTDFILL69_2056 VDD VSS sg13g2_FILL8
XSTDFILL69_2064 VDD VSS sg13g2_FILL8
XSTDFILL69_2072 VDD VSS sg13g2_FILL8
XSTDFILL69_2080 VDD VSS sg13g2_FILL8
XSTDFILL69_2088 VDD VSS sg13g2_FILL8
XSTDFILL69_2096 VDD VSS sg13g2_FILL8
XSTDFILL69_2104 VDD VSS sg13g2_FILL8
XSTDFILL69_2112 VDD VSS sg13g2_FILL8
XSTDFILL69_2120 VDD VSS sg13g2_FILL8
XSTDFILL69_2128 VDD VSS sg13g2_FILL8
XSTDFILL69_2136 VDD VSS sg13g2_FILL8
XSTDFILL69_2144 VDD VSS sg13g2_FILL8
XSTDFILL69_2152 VDD VSS sg13g2_FILL8
XSTDFILL69_2160 VDD VSS sg13g2_FILL8
XSTDFILL69_2168 VDD VSS sg13g2_FILL4
XSTDFILL70_0 VDD VSS sg13g2_FILL8
XSTDFILL70_8 VDD VSS sg13g2_FILL8
XSTDFILL70_16 VDD VSS sg13g2_FILL8
XSTDFILL70_24 VDD VSS sg13g2_FILL8
XSTDFILL70_32 VDD VSS sg13g2_FILL8
XSTDFILL70_40 VDD VSS sg13g2_FILL8
XSTDFILL70_48 VDD VSS sg13g2_FILL8
XSTDFILL70_56 VDD VSS sg13g2_FILL8
XSTDFILL70_64 VDD VSS sg13g2_FILL8
XSTDFILL70_72 VDD VSS sg13g2_FILL8
XSTDFILL70_80 VDD VSS sg13g2_FILL8
XSTDFILL70_88 VDD VSS sg13g2_FILL8
XSTDFILL70_96 VDD VSS sg13g2_FILL8
XSTDFILL70_104 VDD VSS sg13g2_FILL8
XSTDFILL70_112 VDD VSS sg13g2_FILL8
XSTDFILL70_120 VDD VSS sg13g2_FILL8
XSTDFILL70_128 VDD VSS sg13g2_FILL8
XSTDFILL70_136 VDD VSS sg13g2_FILL8
XSTDFILL70_144 VDD VSS sg13g2_FILL8
XSTDFILL70_152 VDD VSS sg13g2_FILL8
XSTDFILL70_160 VDD VSS sg13g2_FILL8
XSTDFILL70_168 VDD VSS sg13g2_FILL8
XSTDFILL70_176 VDD VSS sg13g2_FILL8
XSTDFILL70_184 VDD VSS sg13g2_FILL8
XSTDFILL70_192 VDD VSS sg13g2_FILL8
XSTDFILL70_200 VDD VSS sg13g2_FILL8
XSTDFILL70_208 VDD VSS sg13g2_FILL8
XSTDFILL70_216 VDD VSS sg13g2_FILL8
XSTDFILL70_224 VDD VSS sg13g2_FILL8
XSTDFILL70_232 VDD VSS sg13g2_FILL8
XSTDFILL70_240 VDD VSS sg13g2_FILL8
XSTDFILL70_248 VDD VSS sg13g2_FILL8
XSTDFILL70_256 VDD VSS sg13g2_FILL8
XSTDFILL70_264 VDD VSS sg13g2_FILL8
XSTDFILL70_272 VDD VSS sg13g2_FILL8
XSTDFILL70_280 VDD VSS sg13g2_FILL8
XSTDFILL70_288 VDD VSS sg13g2_FILL8
XSTDFILL70_296 VDD VSS sg13g2_FILL8
XSTDFILL70_304 VDD VSS sg13g2_FILL8
XSTDFILL70_312 VDD VSS sg13g2_FILL8
XSTDFILL70_320 VDD VSS sg13g2_FILL8
XSTDFILL70_328 VDD VSS sg13g2_FILL8
XSTDFILL70_336 VDD VSS sg13g2_FILL8
XSTDFILL70_344 VDD VSS sg13g2_FILL8
XSTDFILL70_352 VDD VSS sg13g2_FILL8
XSTDFILL70_360 VDD VSS sg13g2_FILL8
XSTDFILL70_368 VDD VSS sg13g2_FILL8
XSTDFILL70_376 VDD VSS sg13g2_FILL8
XSTDFILL70_384 VDD VSS sg13g2_FILL8
XSTDFILL70_392 VDD VSS sg13g2_FILL8
XSTDFILL70_400 VDD VSS sg13g2_FILL8
XSTDFILL70_408 VDD VSS sg13g2_FILL8
XSTDFILL70_416 VDD VSS sg13g2_FILL8
XSTDFILL70_424 VDD VSS sg13g2_FILL8
XSTDFILL70_432 VDD VSS sg13g2_FILL8
XSTDFILL70_440 VDD VSS sg13g2_FILL8
XSTDFILL70_448 VDD VSS sg13g2_FILL8
XSTDFILL70_456 VDD VSS sg13g2_FILL8
XSTDFILL70_464 VDD VSS sg13g2_FILL8
XSTDFILL70_472 VDD VSS sg13g2_FILL8
XSTDFILL70_480 VDD VSS sg13g2_FILL8
XSTDFILL70_488 VDD VSS sg13g2_FILL8
XSTDFILL70_496 VDD VSS sg13g2_FILL8
XSTDFILL70_504 VDD VSS sg13g2_FILL8
XSTDFILL70_512 VDD VSS sg13g2_FILL8
XSTDFILL70_520 VDD VSS sg13g2_FILL8
XSTDFILL70_528 VDD VSS sg13g2_FILL8
XSTDFILL70_536 VDD VSS sg13g2_FILL8
XSTDFILL70_544 VDD VSS sg13g2_FILL8
XSTDFILL70_552 VDD VSS sg13g2_FILL8
XSTDFILL70_560 VDD VSS sg13g2_FILL8
XSTDFILL70_568 VDD VSS sg13g2_FILL8
XSTDFILL70_576 VDD VSS sg13g2_FILL8
XSTDFILL70_584 VDD VSS sg13g2_FILL8
XSTDFILL70_592 VDD VSS sg13g2_FILL8
XSTDFILL70_600 VDD VSS sg13g2_FILL8
XSTDFILL70_608 VDD VSS sg13g2_FILL8
XSTDFILL70_616 VDD VSS sg13g2_FILL8
XSTDFILL70_624 VDD VSS sg13g2_FILL8
XSTDFILL70_632 VDD VSS sg13g2_FILL8
XSTDFILL70_640 VDD VSS sg13g2_FILL8
XSTDFILL70_648 VDD VSS sg13g2_FILL8
XSTDFILL70_656 VDD VSS sg13g2_FILL8
XSTDFILL70_664 VDD VSS sg13g2_FILL8
XSTDFILL70_672 VDD VSS sg13g2_FILL8
XSTDFILL70_680 VDD VSS sg13g2_FILL8
XSTDFILL70_688 VDD VSS sg13g2_FILL8
XSTDFILL70_696 VDD VSS sg13g2_FILL8
XSTDFILL70_704 VDD VSS sg13g2_FILL8
XSTDFILL70_712 VDD VSS sg13g2_FILL8
XSTDFILL70_720 VDD VSS sg13g2_FILL8
XSTDFILL70_728 VDD VSS sg13g2_FILL8
XSTDFILL70_736 VDD VSS sg13g2_FILL8
XSTDFILL70_744 VDD VSS sg13g2_FILL8
XSTDFILL70_752 VDD VSS sg13g2_FILL8
XSTDFILL70_760 VDD VSS sg13g2_FILL8
XSTDFILL70_768 VDD VSS sg13g2_FILL8
XSTDFILL70_776 VDD VSS sg13g2_FILL8
XSTDFILL70_784 VDD VSS sg13g2_FILL8
XSTDFILL70_792 VDD VSS sg13g2_FILL8
XSTDFILL70_800 VDD VSS sg13g2_FILL8
XSTDFILL70_808 VDD VSS sg13g2_FILL8
XSTDFILL70_816 VDD VSS sg13g2_FILL8
XSTDFILL70_824 VDD VSS sg13g2_FILL8
XSTDFILL70_832 VDD VSS sg13g2_FILL8
XSTDFILL70_840 VDD VSS sg13g2_FILL8
XSTDFILL70_848 VDD VSS sg13g2_FILL8
XSTDFILL70_856 VDD VSS sg13g2_FILL8
XSTDFILL70_864 VDD VSS sg13g2_FILL8
XSTDFILL70_872 VDD VSS sg13g2_FILL8
XSTDFILL70_880 VDD VSS sg13g2_FILL8
XSTDFILL70_888 VDD VSS sg13g2_FILL8
XSTDFILL70_896 VDD VSS sg13g2_FILL8
XSTDFILL70_904 VDD VSS sg13g2_FILL8
XSTDFILL70_912 VDD VSS sg13g2_FILL8
XSTDFILL70_920 VDD VSS sg13g2_FILL8
XSTDFILL70_928 VDD VSS sg13g2_FILL8
XSTDFILL70_936 VDD VSS sg13g2_FILL8
XSTDFILL70_944 VDD VSS sg13g2_FILL8
XSTDFILL70_952 VDD VSS sg13g2_FILL8
XSTDFILL70_960 VDD VSS sg13g2_FILL8
XSTDFILL70_968 VDD VSS sg13g2_FILL8
XSTDFILL70_976 VDD VSS sg13g2_FILL8
XSTDFILL70_984 VDD VSS sg13g2_FILL8
XSTDFILL70_992 VDD VSS sg13g2_FILL8
XSTDFILL70_1000 VDD VSS sg13g2_FILL8
XSTDFILL70_1008 VDD VSS sg13g2_FILL8
XSTDFILL70_1016 VDD VSS sg13g2_FILL8
XSTDFILL70_1024 VDD VSS sg13g2_FILL8
XSTDFILL70_1032 VDD VSS sg13g2_FILL8
XSTDFILL70_1040 VDD VSS sg13g2_FILL8
XSTDFILL70_1048 VDD VSS sg13g2_FILL8
XSTDFILL70_1056 VDD VSS sg13g2_FILL8
XSTDFILL70_1064 VDD VSS sg13g2_FILL8
XSTDFILL70_1072 VDD VSS sg13g2_FILL8
XSTDFILL70_1080 VDD VSS sg13g2_FILL8
XSTDFILL70_1088 VDD VSS sg13g2_FILL8
XSTDFILL70_1096 VDD VSS sg13g2_FILL8
XSTDFILL70_1104 VDD VSS sg13g2_FILL8
XSTDFILL70_1112 VDD VSS sg13g2_FILL8
XSTDFILL70_1120 VDD VSS sg13g2_FILL8
XSTDFILL70_1128 VDD VSS sg13g2_FILL8
XSTDFILL70_1136 VDD VSS sg13g2_FILL8
XSTDFILL70_1144 VDD VSS sg13g2_FILL8
XSTDFILL70_1152 VDD VSS sg13g2_FILL8
XSTDFILL70_1160 VDD VSS sg13g2_FILL8
XSTDFILL70_1168 VDD VSS sg13g2_FILL8
XSTDFILL70_1176 VDD VSS sg13g2_FILL8
XSTDFILL70_1184 VDD VSS sg13g2_FILL8
XSTDFILL70_1192 VDD VSS sg13g2_FILL8
XSTDFILL70_1200 VDD VSS sg13g2_FILL8
XSTDFILL70_1208 VDD VSS sg13g2_FILL8
XSTDFILL70_1216 VDD VSS sg13g2_FILL8
XSTDFILL70_1224 VDD VSS sg13g2_FILL8
XSTDFILL70_1232 VDD VSS sg13g2_FILL8
XSTDFILL70_1240 VDD VSS sg13g2_FILL8
XSTDFILL70_1248 VDD VSS sg13g2_FILL8
XSTDFILL70_1256 VDD VSS sg13g2_FILL8
XSTDFILL70_1264 VDD VSS sg13g2_FILL8
XSTDFILL70_1272 VDD VSS sg13g2_FILL8
XSTDFILL70_1280 VDD VSS sg13g2_FILL8
XSTDFILL70_1288 VDD VSS sg13g2_FILL8
XSTDFILL70_1296 VDD VSS sg13g2_FILL8
XSTDFILL70_1304 VDD VSS sg13g2_FILL8
XSTDFILL70_1312 VDD VSS sg13g2_FILL8
XSTDFILL70_1320 VDD VSS sg13g2_FILL8
XSTDFILL70_1328 VDD VSS sg13g2_FILL8
XSTDFILL70_1336 VDD VSS sg13g2_FILL8
XSTDFILL70_1344 VDD VSS sg13g2_FILL8
XSTDFILL70_1352 VDD VSS sg13g2_FILL8
XSTDFILL70_1360 VDD VSS sg13g2_FILL8
XSTDFILL70_1368 VDD VSS sg13g2_FILL8
XSTDFILL70_1376 VDD VSS sg13g2_FILL8
XSTDFILL70_1384 VDD VSS sg13g2_FILL8
XSTDFILL70_1392 VDD VSS sg13g2_FILL8
XSTDFILL70_1400 VDD VSS sg13g2_FILL8
XSTDFILL70_1408 VDD VSS sg13g2_FILL8
XSTDFILL70_1416 VDD VSS sg13g2_FILL8
XSTDFILL70_1424 VDD VSS sg13g2_FILL8
XSTDFILL70_1432 VDD VSS sg13g2_FILL8
XSTDFILL70_1440 VDD VSS sg13g2_FILL8
XSTDFILL70_1448 VDD VSS sg13g2_FILL8
XSTDFILL70_1456 VDD VSS sg13g2_FILL8
XSTDFILL70_1464 VDD VSS sg13g2_FILL8
XSTDFILL70_1472 VDD VSS sg13g2_FILL8
XSTDFILL70_1480 VDD VSS sg13g2_FILL8
XSTDFILL70_1488 VDD VSS sg13g2_FILL8
XSTDFILL70_1496 VDD VSS sg13g2_FILL8
XSTDFILL70_1504 VDD VSS sg13g2_FILL8
XSTDFILL70_1512 VDD VSS sg13g2_FILL8
XSTDFILL70_1520 VDD VSS sg13g2_FILL8
XSTDFILL70_1528 VDD VSS sg13g2_FILL8
XSTDFILL70_1536 VDD VSS sg13g2_FILL8
XSTDFILL70_1544 VDD VSS sg13g2_FILL8
XSTDFILL70_1552 VDD VSS sg13g2_FILL8
XSTDFILL70_1560 VDD VSS sg13g2_FILL8
XSTDFILL70_1568 VDD VSS sg13g2_FILL8
XSTDFILL70_1576 VDD VSS sg13g2_FILL8
XSTDFILL70_1584 VDD VSS sg13g2_FILL8
XSTDFILL70_1592 VDD VSS sg13g2_FILL8
XSTDFILL70_1600 VDD VSS sg13g2_FILL8
XSTDFILL70_1608 VDD VSS sg13g2_FILL8
XSTDFILL70_1616 VDD VSS sg13g2_FILL8
XSTDFILL70_1624 VDD VSS sg13g2_FILL8
XSTDFILL70_1632 VDD VSS sg13g2_FILL8
XSTDFILL70_1640 VDD VSS sg13g2_FILL8
XSTDFILL70_1648 VDD VSS sg13g2_FILL8
XSTDFILL70_1656 VDD VSS sg13g2_FILL8
XSTDFILL70_1664 VDD VSS sg13g2_FILL8
XSTDFILL70_1672 VDD VSS sg13g2_FILL8
XSTDFILL70_1680 VDD VSS sg13g2_FILL8
XSTDFILL70_1688 VDD VSS sg13g2_FILL8
XSTDFILL70_1696 VDD VSS sg13g2_FILL8
XSTDFILL70_1704 VDD VSS sg13g2_FILL8
XSTDFILL70_1712 VDD VSS sg13g2_FILL8
XSTDFILL70_1720 VDD VSS sg13g2_FILL8
XSTDFILL70_1728 VDD VSS sg13g2_FILL8
XSTDFILL70_1736 VDD VSS sg13g2_FILL8
XSTDFILL70_1744 VDD VSS sg13g2_FILL8
XSTDFILL70_1752 VDD VSS sg13g2_FILL8
XSTDFILL70_1760 VDD VSS sg13g2_FILL8
XSTDFILL70_1768 VDD VSS sg13g2_FILL8
XSTDFILL70_1776 VDD VSS sg13g2_FILL8
XSTDFILL70_1784 VDD VSS sg13g2_FILL8
XSTDFILL70_1792 VDD VSS sg13g2_FILL8
XSTDFILL70_1800 VDD VSS sg13g2_FILL8
XSTDFILL70_1808 VDD VSS sg13g2_FILL8
XSTDFILL70_1816 VDD VSS sg13g2_FILL8
XSTDFILL70_1824 VDD VSS sg13g2_FILL8
XSTDFILL70_1832 VDD VSS sg13g2_FILL8
XSTDFILL70_1840 VDD VSS sg13g2_FILL8
XSTDFILL70_1848 VDD VSS sg13g2_FILL8
XSTDFILL70_1856 VDD VSS sg13g2_FILL8
XSTDFILL70_1864 VDD VSS sg13g2_FILL8
XSTDFILL70_1872 VDD VSS sg13g2_FILL8
XSTDFILL70_1880 VDD VSS sg13g2_FILL8
XSTDFILL70_1888 VDD VSS sg13g2_FILL8
XSTDFILL70_1896 VDD VSS sg13g2_FILL8
XSTDFILL70_1904 VDD VSS sg13g2_FILL8
XSTDFILL70_1912 VDD VSS sg13g2_FILL8
XSTDFILL70_1920 VDD VSS sg13g2_FILL8
XSTDFILL70_1928 VDD VSS sg13g2_FILL8
XSTDFILL70_1936 VDD VSS sg13g2_FILL8
XSTDFILL70_1944 VDD VSS sg13g2_FILL8
XSTDFILL70_1952 VDD VSS sg13g2_FILL8
XSTDFILL70_1960 VDD VSS sg13g2_FILL8
XSTDFILL70_1968 VDD VSS sg13g2_FILL8
XSTDFILL70_1976 VDD VSS sg13g2_FILL8
XSTDFILL70_1984 VDD VSS sg13g2_FILL8
XSTDFILL70_1992 VDD VSS sg13g2_FILL8
XSTDFILL70_2000 VDD VSS sg13g2_FILL8
XSTDFILL70_2008 VDD VSS sg13g2_FILL8
XSTDFILL70_2016 VDD VSS sg13g2_FILL8
XSTDFILL70_2024 VDD VSS sg13g2_FILL8
XSTDFILL70_2032 VDD VSS sg13g2_FILL8
XSTDFILL70_2040 VDD VSS sg13g2_FILL8
XSTDFILL70_2048 VDD VSS sg13g2_FILL8
XSTDFILL70_2056 VDD VSS sg13g2_FILL8
XSTDFILL70_2064 VDD VSS sg13g2_FILL8
XSTDFILL70_2072 VDD VSS sg13g2_FILL8
XSTDFILL70_2080 VDD VSS sg13g2_FILL8
XSTDFILL70_2088 VDD VSS sg13g2_FILL8
XSTDFILL70_2096 VDD VSS sg13g2_FILL8
XSTDFILL70_2104 VDD VSS sg13g2_FILL8
XSTDFILL70_2112 VDD VSS sg13g2_FILL8
XSTDFILL70_2120 VDD VSS sg13g2_FILL8
XSTDFILL70_2128 VDD VSS sg13g2_FILL8
XSTDFILL70_2136 VDD VSS sg13g2_FILL8
XSTDFILL70_2144 VDD VSS sg13g2_FILL8
XSTDFILL70_2152 VDD VSS sg13g2_FILL8
XSTDFILL70_2160 VDD VSS sg13g2_FILL8
XSTDFILL70_2168 VDD VSS sg13g2_FILL4
XSTDFILL71_0 VDD VSS sg13g2_FILL8
XSTDFILL71_8 VDD VSS sg13g2_FILL8
XSTDFILL71_16 VDD VSS sg13g2_FILL8
XSTDFILL71_24 VDD VSS sg13g2_FILL8
XSTDFILL71_32 VDD VSS sg13g2_FILL8
XSTDFILL71_40 VDD VSS sg13g2_FILL8
XSTDFILL71_48 VDD VSS sg13g2_FILL8
XSTDFILL71_56 VDD VSS sg13g2_FILL8
XSTDFILL71_64 VDD VSS sg13g2_FILL8
XSTDFILL71_72 VDD VSS sg13g2_FILL8
XSTDFILL71_80 VDD VSS sg13g2_FILL8
XSTDFILL71_88 VDD VSS sg13g2_FILL8
XSTDFILL71_96 VDD VSS sg13g2_FILL8
XSTDFILL71_104 VDD VSS sg13g2_FILL8
XSTDFILL71_112 VDD VSS sg13g2_FILL8
XSTDFILL71_120 VDD VSS sg13g2_FILL8
XSTDFILL71_128 VDD VSS sg13g2_FILL8
XSTDFILL71_136 VDD VSS sg13g2_FILL8
XSTDFILL71_144 VDD VSS sg13g2_FILL8
XSTDFILL71_152 VDD VSS sg13g2_FILL8
XSTDFILL71_160 VDD VSS sg13g2_FILL8
XSTDFILL71_168 VDD VSS sg13g2_FILL8
XSTDFILL71_176 VDD VSS sg13g2_FILL8
XSTDFILL71_184 VDD VSS sg13g2_FILL8
XSTDFILL71_192 VDD VSS sg13g2_FILL8
XSTDFILL71_200 VDD VSS sg13g2_FILL8
XSTDFILL71_208 VDD VSS sg13g2_FILL8
XSTDFILL71_216 VDD VSS sg13g2_FILL8
XSTDFILL71_224 VDD VSS sg13g2_FILL8
XSTDFILL71_232 VDD VSS sg13g2_FILL8
XSTDFILL71_240 VDD VSS sg13g2_FILL8
XSTDFILL71_248 VDD VSS sg13g2_FILL8
XSTDFILL71_256 VDD VSS sg13g2_FILL8
XSTDFILL71_264 VDD VSS sg13g2_FILL8
XSTDFILL71_272 VDD VSS sg13g2_FILL8
XSTDFILL71_280 VDD VSS sg13g2_FILL8
XSTDFILL71_288 VDD VSS sg13g2_FILL8
XSTDFILL71_296 VDD VSS sg13g2_FILL8
XSTDFILL71_304 VDD VSS sg13g2_FILL8
XSTDFILL71_312 VDD VSS sg13g2_FILL8
XSTDFILL71_320 VDD VSS sg13g2_FILL8
XSTDFILL71_328 VDD VSS sg13g2_FILL8
XSTDFILL71_336 VDD VSS sg13g2_FILL8
XSTDFILL71_344 VDD VSS sg13g2_FILL8
XSTDFILL71_352 VDD VSS sg13g2_FILL8
XSTDFILL71_360 VDD VSS sg13g2_FILL8
XSTDFILL71_368 VDD VSS sg13g2_FILL8
XSTDFILL71_376 VDD VSS sg13g2_FILL8
XSTDFILL71_384 VDD VSS sg13g2_FILL8
XSTDFILL71_392 VDD VSS sg13g2_FILL8
XSTDFILL71_400 VDD VSS sg13g2_FILL8
XSTDFILL71_408 VDD VSS sg13g2_FILL8
XSTDFILL71_416 VDD VSS sg13g2_FILL8
XSTDFILL71_424 VDD VSS sg13g2_FILL8
XSTDFILL71_432 VDD VSS sg13g2_FILL8
XSTDFILL71_440 VDD VSS sg13g2_FILL8
XSTDFILL71_448 VDD VSS sg13g2_FILL8
XSTDFILL71_456 VDD VSS sg13g2_FILL8
XSTDFILL71_464 VDD VSS sg13g2_FILL8
XSTDFILL71_472 VDD VSS sg13g2_FILL8
XSTDFILL71_480 VDD VSS sg13g2_FILL8
XSTDFILL71_488 VDD VSS sg13g2_FILL8
XSTDFILL71_496 VDD VSS sg13g2_FILL8
XSTDFILL71_504 VDD VSS sg13g2_FILL8
XSTDFILL71_512 VDD VSS sg13g2_FILL8
XSTDFILL71_520 VDD VSS sg13g2_FILL8
XSTDFILL71_528 VDD VSS sg13g2_FILL8
XSTDFILL71_536 VDD VSS sg13g2_FILL8
XSTDFILL71_544 VDD VSS sg13g2_FILL8
XSTDFILL71_552 VDD VSS sg13g2_FILL8
XSTDFILL71_560 VDD VSS sg13g2_FILL8
XSTDFILL71_568 VDD VSS sg13g2_FILL8
XSTDFILL71_576 VDD VSS sg13g2_FILL8
XSTDFILL71_584 VDD VSS sg13g2_FILL8
XSTDFILL71_592 VDD VSS sg13g2_FILL8
XSTDFILL71_600 VDD VSS sg13g2_FILL8
XSTDFILL71_608 VDD VSS sg13g2_FILL8
XSTDFILL71_616 VDD VSS sg13g2_FILL8
XSTDFILL71_624 VDD VSS sg13g2_FILL8
XSTDFILL71_632 VDD VSS sg13g2_FILL8
XSTDFILL71_640 VDD VSS sg13g2_FILL8
XSTDFILL71_648 VDD VSS sg13g2_FILL8
XSTDFILL71_656 VDD VSS sg13g2_FILL8
XSTDFILL71_664 VDD VSS sg13g2_FILL8
XSTDFILL71_672 VDD VSS sg13g2_FILL8
XSTDFILL71_680 VDD VSS sg13g2_FILL8
XSTDFILL71_688 VDD VSS sg13g2_FILL8
XSTDFILL71_696 VDD VSS sg13g2_FILL8
XSTDFILL71_704 VDD VSS sg13g2_FILL8
XSTDFILL71_712 VDD VSS sg13g2_FILL8
XSTDFILL71_720 VDD VSS sg13g2_FILL8
XSTDFILL71_728 VDD VSS sg13g2_FILL8
XSTDFILL71_736 VDD VSS sg13g2_FILL8
XSTDFILL71_744 VDD VSS sg13g2_FILL8
XSTDFILL71_752 VDD VSS sg13g2_FILL8
XSTDFILL71_760 VDD VSS sg13g2_FILL8
XSTDFILL71_768 VDD VSS sg13g2_FILL8
XSTDFILL71_776 VDD VSS sg13g2_FILL8
XSTDFILL71_784 VDD VSS sg13g2_FILL8
XSTDFILL71_792 VDD VSS sg13g2_FILL8
XSTDFILL71_800 VDD VSS sg13g2_FILL8
XSTDFILL71_808 VDD VSS sg13g2_FILL8
XSTDFILL71_816 VDD VSS sg13g2_FILL8
XSTDFILL71_824 VDD VSS sg13g2_FILL8
XSTDFILL71_832 VDD VSS sg13g2_FILL8
XSTDFILL71_840 VDD VSS sg13g2_FILL8
XSTDFILL71_848 VDD VSS sg13g2_FILL8
XSTDFILL71_856 VDD VSS sg13g2_FILL8
XSTDFILL71_864 VDD VSS sg13g2_FILL8
XSTDFILL71_872 VDD VSS sg13g2_FILL8
XSTDFILL71_880 VDD VSS sg13g2_FILL8
XSTDFILL71_888 VDD VSS sg13g2_FILL8
XSTDFILL71_896 VDD VSS sg13g2_FILL8
XSTDFILL71_904 VDD VSS sg13g2_FILL8
XSTDFILL71_912 VDD VSS sg13g2_FILL8
XSTDFILL71_920 VDD VSS sg13g2_FILL8
XSTDFILL71_928 VDD VSS sg13g2_FILL8
XSTDFILL71_936 VDD VSS sg13g2_FILL8
XSTDFILL71_944 VDD VSS sg13g2_FILL8
XSTDFILL71_952 VDD VSS sg13g2_FILL8
XSTDFILL71_960 VDD VSS sg13g2_FILL8
XSTDFILL71_968 VDD VSS sg13g2_FILL8
XSTDFILL71_976 VDD VSS sg13g2_FILL8
XSTDFILL71_984 VDD VSS sg13g2_FILL8
XSTDFILL71_992 VDD VSS sg13g2_FILL8
XSTDFILL71_1000 VDD VSS sg13g2_FILL8
XSTDFILL71_1008 VDD VSS sg13g2_FILL8
XSTDFILL71_1016 VDD VSS sg13g2_FILL8
XSTDFILL71_1024 VDD VSS sg13g2_FILL8
XSTDFILL71_1032 VDD VSS sg13g2_FILL8
XSTDFILL71_1040 VDD VSS sg13g2_FILL8
XSTDFILL71_1048 VDD VSS sg13g2_FILL8
XSTDFILL71_1056 VDD VSS sg13g2_FILL8
XSTDFILL71_1064 VDD VSS sg13g2_FILL8
XSTDFILL71_1072 VDD VSS sg13g2_FILL8
XSTDFILL71_1080 VDD VSS sg13g2_FILL8
XSTDFILL71_1088 VDD VSS sg13g2_FILL8
XSTDFILL71_1096 VDD VSS sg13g2_FILL8
XSTDFILL71_1104 VDD VSS sg13g2_FILL8
XSTDFILL71_1112 VDD VSS sg13g2_FILL8
XSTDFILL71_1120 VDD VSS sg13g2_FILL8
XSTDFILL71_1128 VDD VSS sg13g2_FILL8
XSTDFILL71_1136 VDD VSS sg13g2_FILL8
XSTDFILL71_1144 VDD VSS sg13g2_FILL8
XSTDFILL71_1152 VDD VSS sg13g2_FILL8
XSTDFILL71_1160 VDD VSS sg13g2_FILL8
XSTDFILL71_1168 VDD VSS sg13g2_FILL8
XSTDFILL71_1176 VDD VSS sg13g2_FILL8
XSTDFILL71_1184 VDD VSS sg13g2_FILL8
XSTDFILL71_1192 VDD VSS sg13g2_FILL8
XSTDFILL71_1200 VDD VSS sg13g2_FILL8
XSTDFILL71_1208 VDD VSS sg13g2_FILL8
XSTDFILL71_1216 VDD VSS sg13g2_FILL8
XSTDFILL71_1224 VDD VSS sg13g2_FILL8
XSTDFILL71_1232 VDD VSS sg13g2_FILL8
XSTDFILL71_1240 VDD VSS sg13g2_FILL8
XSTDFILL71_1248 VDD VSS sg13g2_FILL8
XSTDFILL71_1256 VDD VSS sg13g2_FILL8
XSTDFILL71_1264 VDD VSS sg13g2_FILL8
XSTDFILL71_1272 VDD VSS sg13g2_FILL8
XSTDFILL71_1280 VDD VSS sg13g2_FILL8
XSTDFILL71_1288 VDD VSS sg13g2_FILL8
XSTDFILL71_1296 VDD VSS sg13g2_FILL8
XSTDFILL71_1304 VDD VSS sg13g2_FILL8
XSTDFILL71_1312 VDD VSS sg13g2_FILL8
XSTDFILL71_1320 VDD VSS sg13g2_FILL8
XSTDFILL71_1328 VDD VSS sg13g2_FILL8
XSTDFILL71_1336 VDD VSS sg13g2_FILL8
XSTDFILL71_1344 VDD VSS sg13g2_FILL8
XSTDFILL71_1352 VDD VSS sg13g2_FILL8
XSTDFILL71_1360 VDD VSS sg13g2_FILL8
XSTDFILL71_1368 VDD VSS sg13g2_FILL8
XSTDFILL71_1376 VDD VSS sg13g2_FILL8
XSTDFILL71_1384 VDD VSS sg13g2_FILL8
XSTDFILL71_1392 VDD VSS sg13g2_FILL8
XSTDFILL71_1400 VDD VSS sg13g2_FILL8
XSTDFILL71_1408 VDD VSS sg13g2_FILL8
XSTDFILL71_1416 VDD VSS sg13g2_FILL8
XSTDFILL71_1424 VDD VSS sg13g2_FILL8
XSTDFILL71_1432 VDD VSS sg13g2_FILL8
XSTDFILL71_1440 VDD VSS sg13g2_FILL8
XSTDFILL71_1448 VDD VSS sg13g2_FILL8
XSTDFILL71_1456 VDD VSS sg13g2_FILL8
XSTDFILL71_1464 VDD VSS sg13g2_FILL8
XSTDFILL71_1472 VDD VSS sg13g2_FILL8
XSTDFILL71_1480 VDD VSS sg13g2_FILL8
XSTDFILL71_1488 VDD VSS sg13g2_FILL8
XSTDFILL71_1496 VDD VSS sg13g2_FILL8
XSTDFILL71_1504 VDD VSS sg13g2_FILL8
XSTDFILL71_1512 VDD VSS sg13g2_FILL8
XSTDFILL71_1520 VDD VSS sg13g2_FILL8
XSTDFILL71_1528 VDD VSS sg13g2_FILL8
XSTDFILL71_1536 VDD VSS sg13g2_FILL8
XSTDFILL71_1544 VDD VSS sg13g2_FILL8
XSTDFILL71_1552 VDD VSS sg13g2_FILL8
XSTDFILL71_1560 VDD VSS sg13g2_FILL8
XSTDFILL71_1568 VDD VSS sg13g2_FILL8
XSTDFILL71_1576 VDD VSS sg13g2_FILL8
XSTDFILL71_1584 VDD VSS sg13g2_FILL8
XSTDFILL71_1592 VDD VSS sg13g2_FILL8
XSTDFILL71_1600 VDD VSS sg13g2_FILL8
XSTDFILL71_1608 VDD VSS sg13g2_FILL8
XSTDFILL71_1616 VDD VSS sg13g2_FILL8
XSTDFILL71_1624 VDD VSS sg13g2_FILL8
XSTDFILL71_1632 VDD VSS sg13g2_FILL8
XSTDFILL71_1640 VDD VSS sg13g2_FILL8
XSTDFILL71_1648 VDD VSS sg13g2_FILL8
XSTDFILL71_1656 VDD VSS sg13g2_FILL8
XSTDFILL71_1664 VDD VSS sg13g2_FILL8
XSTDFILL71_1672 VDD VSS sg13g2_FILL8
XSTDFILL71_1680 VDD VSS sg13g2_FILL8
XSTDFILL71_1688 VDD VSS sg13g2_FILL8
XSTDFILL71_1696 VDD VSS sg13g2_FILL8
XSTDFILL71_1704 VDD VSS sg13g2_FILL8
XSTDFILL71_1712 VDD VSS sg13g2_FILL8
XSTDFILL71_1720 VDD VSS sg13g2_FILL8
XSTDFILL71_1728 VDD VSS sg13g2_FILL8
XSTDFILL71_1736 VDD VSS sg13g2_FILL8
XSTDFILL71_1744 VDD VSS sg13g2_FILL8
XSTDFILL71_1752 VDD VSS sg13g2_FILL8
XSTDFILL71_1760 VDD VSS sg13g2_FILL8
XSTDFILL71_1768 VDD VSS sg13g2_FILL8
XSTDFILL71_1776 VDD VSS sg13g2_FILL8
XSTDFILL71_1784 VDD VSS sg13g2_FILL8
XSTDFILL71_1792 VDD VSS sg13g2_FILL8
XSTDFILL71_1800 VDD VSS sg13g2_FILL8
XSTDFILL71_1808 VDD VSS sg13g2_FILL8
XSTDFILL71_1816 VDD VSS sg13g2_FILL8
XSTDFILL71_1824 VDD VSS sg13g2_FILL8
XSTDFILL71_1832 VDD VSS sg13g2_FILL8
XSTDFILL71_1840 VDD VSS sg13g2_FILL8
XSTDFILL71_1848 VDD VSS sg13g2_FILL8
XSTDFILL71_1856 VDD VSS sg13g2_FILL8
XSTDFILL71_1864 VDD VSS sg13g2_FILL8
XSTDFILL71_1872 VDD VSS sg13g2_FILL8
XSTDFILL71_1880 VDD VSS sg13g2_FILL8
XSTDFILL71_1888 VDD VSS sg13g2_FILL8
XSTDFILL71_1896 VDD VSS sg13g2_FILL8
XSTDFILL71_1904 VDD VSS sg13g2_FILL8
XSTDFILL71_1912 VDD VSS sg13g2_FILL8
XSTDFILL71_1920 VDD VSS sg13g2_FILL8
XSTDFILL71_1928 VDD VSS sg13g2_FILL8
XSTDFILL71_1936 VDD VSS sg13g2_FILL8
XSTDFILL71_1944 VDD VSS sg13g2_FILL8
XSTDFILL71_1952 VDD VSS sg13g2_FILL8
XSTDFILL71_1960 VDD VSS sg13g2_FILL8
XSTDFILL71_1968 VDD VSS sg13g2_FILL8
XSTDFILL71_1976 VDD VSS sg13g2_FILL8
XSTDFILL71_1984 VDD VSS sg13g2_FILL8
XSTDFILL71_1992 VDD VSS sg13g2_FILL8
XSTDFILL71_2000 VDD VSS sg13g2_FILL8
XSTDFILL71_2008 VDD VSS sg13g2_FILL8
XSTDFILL71_2016 VDD VSS sg13g2_FILL8
XSTDFILL71_2024 VDD VSS sg13g2_FILL8
XSTDFILL71_2032 VDD VSS sg13g2_FILL8
XSTDFILL71_2040 VDD VSS sg13g2_FILL8
XSTDFILL71_2048 VDD VSS sg13g2_FILL8
XSTDFILL71_2056 VDD VSS sg13g2_FILL8
XSTDFILL71_2064 VDD VSS sg13g2_FILL8
XSTDFILL71_2072 VDD VSS sg13g2_FILL8
XSTDFILL71_2080 VDD VSS sg13g2_FILL8
XSTDFILL71_2088 VDD VSS sg13g2_FILL8
XSTDFILL71_2096 VDD VSS sg13g2_FILL8
XSTDFILL71_2104 VDD VSS sg13g2_FILL8
XSTDFILL71_2112 VDD VSS sg13g2_FILL8
XSTDFILL71_2120 VDD VSS sg13g2_FILL8
XSTDFILL71_2128 VDD VSS sg13g2_FILL8
XSTDFILL71_2136 VDD VSS sg13g2_FILL8
XSTDFILL71_2144 VDD VSS sg13g2_FILL8
XSTDFILL71_2152 VDD VSS sg13g2_FILL8
XSTDFILL71_2160 VDD VSS sg13g2_FILL8
XSTDFILL71_2168 VDD VSS sg13g2_FILL4
XSTDFILL72_0 VDD VSS sg13g2_FILL8
XSTDFILL72_8 VDD VSS sg13g2_FILL8
XSTDFILL72_16 VDD VSS sg13g2_FILL8
XSTDFILL72_24 VDD VSS sg13g2_FILL8
XSTDFILL72_32 VDD VSS sg13g2_FILL8
XSTDFILL72_40 VDD VSS sg13g2_FILL8
XSTDFILL72_48 VDD VSS sg13g2_FILL8
XSTDFILL72_56 VDD VSS sg13g2_FILL8
XSTDFILL72_64 VDD VSS sg13g2_FILL8
XSTDFILL72_72 VDD VSS sg13g2_FILL8
XSTDFILL72_80 VDD VSS sg13g2_FILL8
XSTDFILL72_88 VDD VSS sg13g2_FILL8
XSTDFILL72_96 VDD VSS sg13g2_FILL8
XSTDFILL72_104 VDD VSS sg13g2_FILL8
XSTDFILL72_112 VDD VSS sg13g2_FILL8
XSTDFILL72_120 VDD VSS sg13g2_FILL8
XSTDFILL72_128 VDD VSS sg13g2_FILL8
XSTDFILL72_136 VDD VSS sg13g2_FILL8
XSTDFILL72_144 VDD VSS sg13g2_FILL8
XSTDFILL72_152 VDD VSS sg13g2_FILL8
XSTDFILL72_160 VDD VSS sg13g2_FILL8
XSTDFILL72_168 VDD VSS sg13g2_FILL8
XSTDFILL72_176 VDD VSS sg13g2_FILL8
XSTDFILL72_184 VDD VSS sg13g2_FILL8
XSTDFILL72_192 VDD VSS sg13g2_FILL8
XSTDFILL72_200 VDD VSS sg13g2_FILL8
XSTDFILL72_208 VDD VSS sg13g2_FILL8
XSTDFILL72_216 VDD VSS sg13g2_FILL8
XSTDFILL72_224 VDD VSS sg13g2_FILL8
XSTDFILL72_232 VDD VSS sg13g2_FILL8
XSTDFILL72_240 VDD VSS sg13g2_FILL8
XSTDFILL72_248 VDD VSS sg13g2_FILL8
XSTDFILL72_256 VDD VSS sg13g2_FILL8
XSTDFILL72_264 VDD VSS sg13g2_FILL8
XSTDFILL72_272 VDD VSS sg13g2_FILL8
XSTDFILL72_280 VDD VSS sg13g2_FILL8
XSTDFILL72_288 VDD VSS sg13g2_FILL8
XSTDFILL72_296 VDD VSS sg13g2_FILL8
XSTDFILL72_304 VDD VSS sg13g2_FILL8
XSTDFILL72_312 VDD VSS sg13g2_FILL8
XSTDFILL72_320 VDD VSS sg13g2_FILL8
XSTDFILL72_328 VDD VSS sg13g2_FILL8
XSTDFILL72_336 VDD VSS sg13g2_FILL8
XSTDFILL72_344 VDD VSS sg13g2_FILL8
XSTDFILL72_352 VDD VSS sg13g2_FILL8
XSTDFILL72_360 VDD VSS sg13g2_FILL8
XSTDFILL72_368 VDD VSS sg13g2_FILL8
XSTDFILL72_376 VDD VSS sg13g2_FILL8
XSTDFILL72_384 VDD VSS sg13g2_FILL8
XSTDFILL72_392 VDD VSS sg13g2_FILL8
XSTDFILL72_400 VDD VSS sg13g2_FILL8
XSTDFILL72_408 VDD VSS sg13g2_FILL8
XSTDFILL72_416 VDD VSS sg13g2_FILL8
XSTDFILL72_424 VDD VSS sg13g2_FILL8
XSTDFILL72_432 VDD VSS sg13g2_FILL8
XSTDFILL72_440 VDD VSS sg13g2_FILL8
XSTDFILL72_448 VDD VSS sg13g2_FILL8
XSTDFILL72_456 VDD VSS sg13g2_FILL8
XSTDFILL72_464 VDD VSS sg13g2_FILL8
XSTDFILL72_472 VDD VSS sg13g2_FILL8
XSTDFILL72_480 VDD VSS sg13g2_FILL8
XSTDFILL72_488 VDD VSS sg13g2_FILL8
XSTDFILL72_496 VDD VSS sg13g2_FILL8
XSTDFILL72_504 VDD VSS sg13g2_FILL8
XSTDFILL72_512 VDD VSS sg13g2_FILL8
XSTDFILL72_520 VDD VSS sg13g2_FILL8
XSTDFILL72_528 VDD VSS sg13g2_FILL8
XSTDFILL72_536 VDD VSS sg13g2_FILL8
XSTDFILL72_544 VDD VSS sg13g2_FILL8
XSTDFILL72_552 VDD VSS sg13g2_FILL8
XSTDFILL72_560 VDD VSS sg13g2_FILL8
XSTDFILL72_568 VDD VSS sg13g2_FILL8
XSTDFILL72_576 VDD VSS sg13g2_FILL8
XSTDFILL72_584 VDD VSS sg13g2_FILL8
XSTDFILL72_592 VDD VSS sg13g2_FILL8
XSTDFILL72_600 VDD VSS sg13g2_FILL8
XSTDFILL72_608 VDD VSS sg13g2_FILL8
XSTDFILL72_616 VDD VSS sg13g2_FILL8
XSTDFILL72_624 VDD VSS sg13g2_FILL8
XSTDFILL72_632 VDD VSS sg13g2_FILL8
XSTDFILL72_640 VDD VSS sg13g2_FILL8
XSTDFILL72_648 VDD VSS sg13g2_FILL8
XSTDFILL72_656 VDD VSS sg13g2_FILL8
XSTDFILL72_664 VDD VSS sg13g2_FILL8
XSTDFILL72_672 VDD VSS sg13g2_FILL8
XSTDFILL72_680 VDD VSS sg13g2_FILL8
XSTDFILL72_688 VDD VSS sg13g2_FILL8
XSTDFILL72_696 VDD VSS sg13g2_FILL8
XSTDFILL72_704 VDD VSS sg13g2_FILL8
XSTDFILL72_712 VDD VSS sg13g2_FILL8
XSTDFILL72_720 VDD VSS sg13g2_FILL8
XSTDFILL72_728 VDD VSS sg13g2_FILL8
XSTDFILL72_736 VDD VSS sg13g2_FILL8
XSTDFILL72_744 VDD VSS sg13g2_FILL8
XSTDFILL72_752 VDD VSS sg13g2_FILL8
XSTDFILL72_760 VDD VSS sg13g2_FILL8
XSTDFILL72_768 VDD VSS sg13g2_FILL8
XSTDFILL72_776 VDD VSS sg13g2_FILL8
XSTDFILL72_784 VDD VSS sg13g2_FILL8
XSTDFILL72_792 VDD VSS sg13g2_FILL8
XSTDFILL72_800 VDD VSS sg13g2_FILL8
XSTDFILL72_808 VDD VSS sg13g2_FILL8
XSTDFILL72_816 VDD VSS sg13g2_FILL8
XSTDFILL72_824 VDD VSS sg13g2_FILL8
XSTDFILL72_832 VDD VSS sg13g2_FILL8
XSTDFILL72_840 VDD VSS sg13g2_FILL8
XSTDFILL72_848 VDD VSS sg13g2_FILL8
XSTDFILL72_856 VDD VSS sg13g2_FILL8
XSTDFILL72_864 VDD VSS sg13g2_FILL8
XSTDFILL72_872 VDD VSS sg13g2_FILL8
XSTDFILL72_880 VDD VSS sg13g2_FILL8
XSTDFILL72_888 VDD VSS sg13g2_FILL8
XSTDFILL72_896 VDD VSS sg13g2_FILL8
XSTDFILL72_904 VDD VSS sg13g2_FILL8
XSTDFILL72_912 VDD VSS sg13g2_FILL8
XSTDFILL72_920 VDD VSS sg13g2_FILL8
XSTDFILL72_928 VDD VSS sg13g2_FILL8
XSTDFILL72_936 VDD VSS sg13g2_FILL8
XSTDFILL72_944 VDD VSS sg13g2_FILL8
XSTDFILL72_952 VDD VSS sg13g2_FILL8
XSTDFILL72_960 VDD VSS sg13g2_FILL8
XSTDFILL72_968 VDD VSS sg13g2_FILL8
XSTDFILL72_976 VDD VSS sg13g2_FILL8
XSTDFILL72_984 VDD VSS sg13g2_FILL8
XSTDFILL72_992 VDD VSS sg13g2_FILL8
XSTDFILL72_1000 VDD VSS sg13g2_FILL8
XSTDFILL72_1008 VDD VSS sg13g2_FILL8
XSTDFILL72_1016 VDD VSS sg13g2_FILL8
XSTDFILL72_1024 VDD VSS sg13g2_FILL8
XSTDFILL72_1032 VDD VSS sg13g2_FILL8
XSTDFILL72_1040 VDD VSS sg13g2_FILL8
XSTDFILL72_1048 VDD VSS sg13g2_FILL8
XSTDFILL72_1056 VDD VSS sg13g2_FILL8
XSTDFILL72_1064 VDD VSS sg13g2_FILL8
XSTDFILL72_1072 VDD VSS sg13g2_FILL8
XSTDFILL72_1080 VDD VSS sg13g2_FILL8
XSTDFILL72_1088 VDD VSS sg13g2_FILL8
XSTDFILL72_1096 VDD VSS sg13g2_FILL8
XSTDFILL72_1104 VDD VSS sg13g2_FILL8
XSTDFILL72_1112 VDD VSS sg13g2_FILL8
XSTDFILL72_1120 VDD VSS sg13g2_FILL8
XSTDFILL72_1128 VDD VSS sg13g2_FILL8
XSTDFILL72_1136 VDD VSS sg13g2_FILL8
XSTDFILL72_1144 VDD VSS sg13g2_FILL8
XSTDFILL72_1152 VDD VSS sg13g2_FILL8
XSTDFILL72_1160 VDD VSS sg13g2_FILL8
XSTDFILL72_1168 VDD VSS sg13g2_FILL8
XSTDFILL72_1176 VDD VSS sg13g2_FILL8
XSTDFILL72_1184 VDD VSS sg13g2_FILL8
XSTDFILL72_1192 VDD VSS sg13g2_FILL8
XSTDFILL72_1200 VDD VSS sg13g2_FILL8
XSTDFILL72_1208 VDD VSS sg13g2_FILL8
XSTDFILL72_1216 VDD VSS sg13g2_FILL8
XSTDFILL72_1224 VDD VSS sg13g2_FILL8
XSTDFILL72_1232 VDD VSS sg13g2_FILL8
XSTDFILL72_1240 VDD VSS sg13g2_FILL8
XSTDFILL72_1248 VDD VSS sg13g2_FILL8
XSTDFILL72_1256 VDD VSS sg13g2_FILL8
XSTDFILL72_1264 VDD VSS sg13g2_FILL8
XSTDFILL72_1272 VDD VSS sg13g2_FILL8
XSTDFILL72_1280 VDD VSS sg13g2_FILL8
XSTDFILL72_1288 VDD VSS sg13g2_FILL8
XSTDFILL72_1296 VDD VSS sg13g2_FILL8
XSTDFILL72_1304 VDD VSS sg13g2_FILL8
XSTDFILL72_1312 VDD VSS sg13g2_FILL8
XSTDFILL72_1320 VDD VSS sg13g2_FILL8
XSTDFILL72_1328 VDD VSS sg13g2_FILL8
XSTDFILL72_1336 VDD VSS sg13g2_FILL8
XSTDFILL72_1344 VDD VSS sg13g2_FILL8
XSTDFILL72_1352 VDD VSS sg13g2_FILL8
XSTDFILL72_1360 VDD VSS sg13g2_FILL8
XSTDFILL72_1368 VDD VSS sg13g2_FILL8
XSTDFILL72_1376 VDD VSS sg13g2_FILL8
XSTDFILL72_1384 VDD VSS sg13g2_FILL8
XSTDFILL72_1392 VDD VSS sg13g2_FILL8
XSTDFILL72_1400 VDD VSS sg13g2_FILL8
XSTDFILL72_1408 VDD VSS sg13g2_FILL8
XSTDFILL72_1416 VDD VSS sg13g2_FILL8
XSTDFILL72_1424 VDD VSS sg13g2_FILL8
XSTDFILL72_1432 VDD VSS sg13g2_FILL8
XSTDFILL72_1440 VDD VSS sg13g2_FILL8
XSTDFILL72_1448 VDD VSS sg13g2_FILL8
XSTDFILL72_1456 VDD VSS sg13g2_FILL8
XSTDFILL72_1464 VDD VSS sg13g2_FILL8
XSTDFILL72_1472 VDD VSS sg13g2_FILL8
XSTDFILL72_1480 VDD VSS sg13g2_FILL8
XSTDFILL72_1488 VDD VSS sg13g2_FILL8
XSTDFILL72_1496 VDD VSS sg13g2_FILL8
XSTDFILL72_1504 VDD VSS sg13g2_FILL8
XSTDFILL72_1512 VDD VSS sg13g2_FILL8
XSTDFILL72_1520 VDD VSS sg13g2_FILL8
XSTDFILL72_1528 VDD VSS sg13g2_FILL8
XSTDFILL72_1536 VDD VSS sg13g2_FILL8
XSTDFILL72_1544 VDD VSS sg13g2_FILL8
XSTDFILL72_1552 VDD VSS sg13g2_FILL8
XSTDFILL72_1560 VDD VSS sg13g2_FILL8
XSTDFILL72_1568 VDD VSS sg13g2_FILL8
XSTDFILL72_1576 VDD VSS sg13g2_FILL8
XSTDFILL72_1584 VDD VSS sg13g2_FILL8
XSTDFILL72_1592 VDD VSS sg13g2_FILL8
XSTDFILL72_1600 VDD VSS sg13g2_FILL8
XSTDFILL72_1608 VDD VSS sg13g2_FILL8
XSTDFILL72_1616 VDD VSS sg13g2_FILL8
XSTDFILL72_1624 VDD VSS sg13g2_FILL8
XSTDFILL72_1632 VDD VSS sg13g2_FILL8
XSTDFILL72_1640 VDD VSS sg13g2_FILL8
XSTDFILL72_1648 VDD VSS sg13g2_FILL8
XSTDFILL72_1656 VDD VSS sg13g2_FILL8
XSTDFILL72_1664 VDD VSS sg13g2_FILL8
XSTDFILL72_1672 VDD VSS sg13g2_FILL8
XSTDFILL72_1680 VDD VSS sg13g2_FILL8
XSTDFILL72_1688 VDD VSS sg13g2_FILL8
XSTDFILL72_1696 VDD VSS sg13g2_FILL8
XSTDFILL72_1704 VDD VSS sg13g2_FILL8
XSTDFILL72_1712 VDD VSS sg13g2_FILL8
XSTDFILL72_1720 VDD VSS sg13g2_FILL8
XSTDFILL72_1728 VDD VSS sg13g2_FILL8
XSTDFILL72_1736 VDD VSS sg13g2_FILL8
XSTDFILL72_1744 VDD VSS sg13g2_FILL8
XSTDFILL72_1752 VDD VSS sg13g2_FILL8
XSTDFILL72_1760 VDD VSS sg13g2_FILL8
XSTDFILL72_1768 VDD VSS sg13g2_FILL8
XSTDFILL72_1776 VDD VSS sg13g2_FILL8
XSTDFILL72_1784 VDD VSS sg13g2_FILL8
XSTDFILL72_1792 VDD VSS sg13g2_FILL8
XSTDFILL72_1800 VDD VSS sg13g2_FILL8
XSTDFILL72_1808 VDD VSS sg13g2_FILL8
XSTDFILL72_1816 VDD VSS sg13g2_FILL8
XSTDFILL72_1824 VDD VSS sg13g2_FILL8
XSTDFILL72_1832 VDD VSS sg13g2_FILL8
XSTDFILL72_1840 VDD VSS sg13g2_FILL8
XSTDFILL72_1848 VDD VSS sg13g2_FILL8
XSTDFILL72_1856 VDD VSS sg13g2_FILL8
XSTDFILL72_1864 VDD VSS sg13g2_FILL8
XSTDFILL72_1872 VDD VSS sg13g2_FILL8
XSTDFILL72_1880 VDD VSS sg13g2_FILL8
XSTDFILL72_1888 VDD VSS sg13g2_FILL8
XSTDFILL72_1896 VDD VSS sg13g2_FILL8
XSTDFILL72_1904 VDD VSS sg13g2_FILL8
XSTDFILL72_1912 VDD VSS sg13g2_FILL8
XSTDFILL72_1920 VDD VSS sg13g2_FILL8
XSTDFILL72_1928 VDD VSS sg13g2_FILL8
XSTDFILL72_1936 VDD VSS sg13g2_FILL8
XSTDFILL72_1944 VDD VSS sg13g2_FILL8
XSTDFILL72_1952 VDD VSS sg13g2_FILL8
XSTDFILL72_1960 VDD VSS sg13g2_FILL8
XSTDFILL72_1968 VDD VSS sg13g2_FILL8
XSTDFILL72_1976 VDD VSS sg13g2_FILL8
XSTDFILL72_1984 VDD VSS sg13g2_FILL8
XSTDFILL72_1992 VDD VSS sg13g2_FILL8
XSTDFILL72_2000 VDD VSS sg13g2_FILL8
XSTDFILL72_2008 VDD VSS sg13g2_FILL8
XSTDFILL72_2016 VDD VSS sg13g2_FILL8
XSTDFILL72_2024 VDD VSS sg13g2_FILL8
XSTDFILL72_2032 VDD VSS sg13g2_FILL8
XSTDFILL72_2040 VDD VSS sg13g2_FILL8
XSTDFILL72_2048 VDD VSS sg13g2_FILL8
XSTDFILL72_2056 VDD VSS sg13g2_FILL8
XSTDFILL72_2064 VDD VSS sg13g2_FILL8
XSTDFILL72_2072 VDD VSS sg13g2_FILL8
XSTDFILL72_2080 VDD VSS sg13g2_FILL8
XSTDFILL72_2088 VDD VSS sg13g2_FILL8
XSTDFILL72_2096 VDD VSS sg13g2_FILL8
XSTDFILL72_2104 VDD VSS sg13g2_FILL8
XSTDFILL72_2112 VDD VSS sg13g2_FILL8
XSTDFILL72_2120 VDD VSS sg13g2_FILL8
XSTDFILL72_2128 VDD VSS sg13g2_FILL8
XSTDFILL72_2136 VDD VSS sg13g2_FILL8
XSTDFILL72_2144 VDD VSS sg13g2_FILL8
XSTDFILL72_2152 VDD VSS sg13g2_FILL8
XSTDFILL72_2160 VDD VSS sg13g2_FILL8
XSTDFILL72_2168 VDD VSS sg13g2_FILL4
XSTDFILL73_0 VDD VSS sg13g2_FILL8
XSTDFILL73_8 VDD VSS sg13g2_FILL8
XSTDFILL73_16 VDD VSS sg13g2_FILL8
XSTDFILL73_24 VDD VSS sg13g2_FILL8
XSTDFILL73_32 VDD VSS sg13g2_FILL8
XSTDFILL73_40 VDD VSS sg13g2_FILL8
XSTDFILL73_48 VDD VSS sg13g2_FILL8
XSTDFILL73_56 VDD VSS sg13g2_FILL8
XSTDFILL73_64 VDD VSS sg13g2_FILL8
XSTDFILL73_72 VDD VSS sg13g2_FILL8
XSTDFILL73_80 VDD VSS sg13g2_FILL8
XSTDFILL73_88 VDD VSS sg13g2_FILL8
XSTDFILL73_96 VDD VSS sg13g2_FILL8
XSTDFILL73_104 VDD VSS sg13g2_FILL8
XSTDFILL73_112 VDD VSS sg13g2_FILL8
XSTDFILL73_120 VDD VSS sg13g2_FILL8
XSTDFILL73_128 VDD VSS sg13g2_FILL8
XSTDFILL73_136 VDD VSS sg13g2_FILL8
XSTDFILL73_144 VDD VSS sg13g2_FILL8
XSTDFILL73_152 VDD VSS sg13g2_FILL8
XSTDFILL73_160 VDD VSS sg13g2_FILL8
XSTDFILL73_168 VDD VSS sg13g2_FILL8
XSTDFILL73_176 VDD VSS sg13g2_FILL8
XSTDFILL73_184 VDD VSS sg13g2_FILL8
XSTDFILL73_192 VDD VSS sg13g2_FILL8
XSTDFILL73_200 VDD VSS sg13g2_FILL8
XSTDFILL73_208 VDD VSS sg13g2_FILL8
XSTDFILL73_216 VDD VSS sg13g2_FILL8
XSTDFILL73_224 VDD VSS sg13g2_FILL8
XSTDFILL73_232 VDD VSS sg13g2_FILL8
XSTDFILL73_240 VDD VSS sg13g2_FILL8
XSTDFILL73_248 VDD VSS sg13g2_FILL8
XSTDFILL73_256 VDD VSS sg13g2_FILL8
XSTDFILL73_264 VDD VSS sg13g2_FILL8
XSTDFILL73_272 VDD VSS sg13g2_FILL8
XSTDFILL73_280 VDD VSS sg13g2_FILL8
XSTDFILL73_288 VDD VSS sg13g2_FILL8
XSTDFILL73_296 VDD VSS sg13g2_FILL8
XSTDFILL73_304 VDD VSS sg13g2_FILL8
XSTDFILL73_312 VDD VSS sg13g2_FILL8
XSTDFILL73_320 VDD VSS sg13g2_FILL8
XSTDFILL73_328 VDD VSS sg13g2_FILL8
XSTDFILL73_336 VDD VSS sg13g2_FILL8
XSTDFILL73_344 VDD VSS sg13g2_FILL8
XSTDFILL73_352 VDD VSS sg13g2_FILL8
XSTDFILL73_360 VDD VSS sg13g2_FILL8
XSTDFILL73_368 VDD VSS sg13g2_FILL8
XSTDFILL73_376 VDD VSS sg13g2_FILL8
XSTDFILL73_384 VDD VSS sg13g2_FILL8
XSTDFILL73_392 VDD VSS sg13g2_FILL8
XSTDFILL73_400 VDD VSS sg13g2_FILL8
XSTDFILL73_408 VDD VSS sg13g2_FILL8
XSTDFILL73_416 VDD VSS sg13g2_FILL8
XSTDFILL73_424 VDD VSS sg13g2_FILL8
XSTDFILL73_432 VDD VSS sg13g2_FILL8
XSTDFILL73_440 VDD VSS sg13g2_FILL8
XSTDFILL73_448 VDD VSS sg13g2_FILL8
XSTDFILL73_456 VDD VSS sg13g2_FILL8
XSTDFILL73_464 VDD VSS sg13g2_FILL8
XSTDFILL73_472 VDD VSS sg13g2_FILL8
XSTDFILL73_480 VDD VSS sg13g2_FILL8
XSTDFILL73_488 VDD VSS sg13g2_FILL8
XSTDFILL73_496 VDD VSS sg13g2_FILL8
XSTDFILL73_504 VDD VSS sg13g2_FILL8
XSTDFILL73_512 VDD VSS sg13g2_FILL8
XSTDFILL73_520 VDD VSS sg13g2_FILL8
XSTDFILL73_528 VDD VSS sg13g2_FILL8
XSTDFILL73_536 VDD VSS sg13g2_FILL8
XSTDFILL73_544 VDD VSS sg13g2_FILL8
XSTDFILL73_552 VDD VSS sg13g2_FILL8
XSTDFILL73_560 VDD VSS sg13g2_FILL8
XSTDFILL73_568 VDD VSS sg13g2_FILL8
XSTDFILL73_576 VDD VSS sg13g2_FILL8
XSTDFILL73_584 VDD VSS sg13g2_FILL8
XSTDFILL73_592 VDD VSS sg13g2_FILL8
XSTDFILL73_600 VDD VSS sg13g2_FILL8
XSTDFILL73_608 VDD VSS sg13g2_FILL8
XSTDFILL73_616 VDD VSS sg13g2_FILL8
XSTDFILL73_624 VDD VSS sg13g2_FILL8
XSTDFILL73_632 VDD VSS sg13g2_FILL8
XSTDFILL73_640 VDD VSS sg13g2_FILL8
XSTDFILL73_648 VDD VSS sg13g2_FILL8
XSTDFILL73_656 VDD VSS sg13g2_FILL8
XSTDFILL73_664 VDD VSS sg13g2_FILL8
XSTDFILL73_672 VDD VSS sg13g2_FILL8
XSTDFILL73_680 VDD VSS sg13g2_FILL8
XSTDFILL73_688 VDD VSS sg13g2_FILL8
XSTDFILL73_696 VDD VSS sg13g2_FILL8
XSTDFILL73_704 VDD VSS sg13g2_FILL8
XSTDFILL73_712 VDD VSS sg13g2_FILL8
XSTDFILL73_720 VDD VSS sg13g2_FILL8
XSTDFILL73_728 VDD VSS sg13g2_FILL8
XSTDFILL73_736 VDD VSS sg13g2_FILL8
XSTDFILL73_744 VDD VSS sg13g2_FILL8
XSTDFILL73_752 VDD VSS sg13g2_FILL8
XSTDFILL73_760 VDD VSS sg13g2_FILL8
XSTDFILL73_768 VDD VSS sg13g2_FILL8
XSTDFILL73_776 VDD VSS sg13g2_FILL8
XSTDFILL73_784 VDD VSS sg13g2_FILL8
XSTDFILL73_792 VDD VSS sg13g2_FILL8
XSTDFILL73_800 VDD VSS sg13g2_FILL8
XSTDFILL73_808 VDD VSS sg13g2_FILL8
XSTDFILL73_816 VDD VSS sg13g2_FILL8
XSTDFILL73_824 VDD VSS sg13g2_FILL8
XSTDFILL73_832 VDD VSS sg13g2_FILL8
XSTDFILL73_840 VDD VSS sg13g2_FILL8
XSTDFILL73_848 VDD VSS sg13g2_FILL8
XSTDFILL73_856 VDD VSS sg13g2_FILL8
XSTDFILL73_864 VDD VSS sg13g2_FILL8
XSTDFILL73_872 VDD VSS sg13g2_FILL8
XSTDFILL73_880 VDD VSS sg13g2_FILL8
XSTDFILL73_888 VDD VSS sg13g2_FILL8
XSTDFILL73_896 VDD VSS sg13g2_FILL8
XSTDFILL73_904 VDD VSS sg13g2_FILL8
XSTDFILL73_912 VDD VSS sg13g2_FILL8
XSTDFILL73_920 VDD VSS sg13g2_FILL8
XSTDFILL73_928 VDD VSS sg13g2_FILL8
XSTDFILL73_936 VDD VSS sg13g2_FILL8
XSTDFILL73_944 VDD VSS sg13g2_FILL8
XSTDFILL73_952 VDD VSS sg13g2_FILL8
XSTDFILL73_960 VDD VSS sg13g2_FILL8
XSTDFILL73_968 VDD VSS sg13g2_FILL8
XSTDFILL73_976 VDD VSS sg13g2_FILL8
XSTDFILL73_984 VDD VSS sg13g2_FILL8
XSTDFILL73_992 VDD VSS sg13g2_FILL8
XSTDFILL73_1000 VDD VSS sg13g2_FILL8
XSTDFILL73_1008 VDD VSS sg13g2_FILL8
XSTDFILL73_1016 VDD VSS sg13g2_FILL8
XSTDFILL73_1024 VDD VSS sg13g2_FILL8
XSTDFILL73_1032 VDD VSS sg13g2_FILL8
XSTDFILL73_1040 VDD VSS sg13g2_FILL8
XSTDFILL73_1048 VDD VSS sg13g2_FILL8
XSTDFILL73_1056 VDD VSS sg13g2_FILL8
XSTDFILL73_1064 VDD VSS sg13g2_FILL8
XSTDFILL73_1072 VDD VSS sg13g2_FILL8
XSTDFILL73_1080 VDD VSS sg13g2_FILL8
XSTDFILL73_1088 VDD VSS sg13g2_FILL8
XSTDFILL73_1096 VDD VSS sg13g2_FILL8
XSTDFILL73_1104 VDD VSS sg13g2_FILL8
XSTDFILL73_1112 VDD VSS sg13g2_FILL8
XSTDFILL73_1120 VDD VSS sg13g2_FILL8
XSTDFILL73_1128 VDD VSS sg13g2_FILL8
XSTDFILL73_1136 VDD VSS sg13g2_FILL8
XSTDFILL73_1144 VDD VSS sg13g2_FILL8
XSTDFILL73_1152 VDD VSS sg13g2_FILL8
XSTDFILL73_1160 VDD VSS sg13g2_FILL8
XSTDFILL73_1168 VDD VSS sg13g2_FILL8
XSTDFILL73_1176 VDD VSS sg13g2_FILL8
XSTDFILL73_1184 VDD VSS sg13g2_FILL8
XSTDFILL73_1192 VDD VSS sg13g2_FILL8
XSTDFILL73_1200 VDD VSS sg13g2_FILL8
XSTDFILL73_1208 VDD VSS sg13g2_FILL8
XSTDFILL73_1216 VDD VSS sg13g2_FILL8
XSTDFILL73_1224 VDD VSS sg13g2_FILL8
XSTDFILL73_1232 VDD VSS sg13g2_FILL8
XSTDFILL73_1240 VDD VSS sg13g2_FILL8
XSTDFILL73_1248 VDD VSS sg13g2_FILL8
XSTDFILL73_1256 VDD VSS sg13g2_FILL8
XSTDFILL73_1264 VDD VSS sg13g2_FILL8
XSTDFILL73_1272 VDD VSS sg13g2_FILL8
XSTDFILL73_1280 VDD VSS sg13g2_FILL8
XSTDFILL73_1288 VDD VSS sg13g2_FILL8
XSTDFILL73_1296 VDD VSS sg13g2_FILL8
XSTDFILL73_1304 VDD VSS sg13g2_FILL8
XSTDFILL73_1312 VDD VSS sg13g2_FILL8
XSTDFILL73_1320 VDD VSS sg13g2_FILL8
XSTDFILL73_1328 VDD VSS sg13g2_FILL8
XSTDFILL73_1336 VDD VSS sg13g2_FILL8
XSTDFILL73_1344 VDD VSS sg13g2_FILL8
XSTDFILL73_1352 VDD VSS sg13g2_FILL8
XSTDFILL73_1360 VDD VSS sg13g2_FILL8
XSTDFILL73_1368 VDD VSS sg13g2_FILL8
XSTDFILL73_1376 VDD VSS sg13g2_FILL8
XSTDFILL73_1384 VDD VSS sg13g2_FILL8
XSTDFILL73_1392 VDD VSS sg13g2_FILL8
XSTDFILL73_1400 VDD VSS sg13g2_FILL8
XSTDFILL73_1408 VDD VSS sg13g2_FILL8
XSTDFILL73_1416 VDD VSS sg13g2_FILL8
XSTDFILL73_1424 VDD VSS sg13g2_FILL8
XSTDFILL73_1432 VDD VSS sg13g2_FILL8
XSTDFILL73_1440 VDD VSS sg13g2_FILL8
XSTDFILL73_1448 VDD VSS sg13g2_FILL8
XSTDFILL73_1456 VDD VSS sg13g2_FILL8
XSTDFILL73_1464 VDD VSS sg13g2_FILL8
XSTDFILL73_1472 VDD VSS sg13g2_FILL8
XSTDFILL73_1480 VDD VSS sg13g2_FILL8
XSTDFILL73_1488 VDD VSS sg13g2_FILL8
XSTDFILL73_1496 VDD VSS sg13g2_FILL8
XSTDFILL73_1504 VDD VSS sg13g2_FILL8
XSTDFILL73_1512 VDD VSS sg13g2_FILL8
XSTDFILL73_1520 VDD VSS sg13g2_FILL8
XSTDFILL73_1528 VDD VSS sg13g2_FILL8
XSTDFILL73_1536 VDD VSS sg13g2_FILL8
XSTDFILL73_1544 VDD VSS sg13g2_FILL8
XSTDFILL73_1552 VDD VSS sg13g2_FILL8
XSTDFILL73_1560 VDD VSS sg13g2_FILL8
XSTDFILL73_1568 VDD VSS sg13g2_FILL8
XSTDFILL73_1576 VDD VSS sg13g2_FILL8
XSTDFILL73_1584 VDD VSS sg13g2_FILL8
XSTDFILL73_1592 VDD VSS sg13g2_FILL8
XSTDFILL73_1600 VDD VSS sg13g2_FILL8
XSTDFILL73_1608 VDD VSS sg13g2_FILL8
XSTDFILL73_1616 VDD VSS sg13g2_FILL8
XSTDFILL73_1624 VDD VSS sg13g2_FILL8
XSTDFILL73_1632 VDD VSS sg13g2_FILL8
XSTDFILL73_1640 VDD VSS sg13g2_FILL8
XSTDFILL73_1648 VDD VSS sg13g2_FILL8
XSTDFILL73_1656 VDD VSS sg13g2_FILL8
XSTDFILL73_1664 VDD VSS sg13g2_FILL8
XSTDFILL73_1672 VDD VSS sg13g2_FILL8
XSTDFILL73_1680 VDD VSS sg13g2_FILL8
XSTDFILL73_1688 VDD VSS sg13g2_FILL8
XSTDFILL73_1696 VDD VSS sg13g2_FILL8
XSTDFILL73_1704 VDD VSS sg13g2_FILL8
XSTDFILL73_1712 VDD VSS sg13g2_FILL8
XSTDFILL73_1720 VDD VSS sg13g2_FILL8
XSTDFILL73_1728 VDD VSS sg13g2_FILL8
XSTDFILL73_1736 VDD VSS sg13g2_FILL8
XSTDFILL73_1744 VDD VSS sg13g2_FILL8
XSTDFILL73_1752 VDD VSS sg13g2_FILL8
XSTDFILL73_1760 VDD VSS sg13g2_FILL8
XSTDFILL73_1768 VDD VSS sg13g2_FILL8
XSTDFILL73_1776 VDD VSS sg13g2_FILL8
XSTDFILL73_1784 VDD VSS sg13g2_FILL8
XSTDFILL73_1792 VDD VSS sg13g2_FILL8
XSTDFILL73_1800 VDD VSS sg13g2_FILL8
XSTDFILL73_1808 VDD VSS sg13g2_FILL8
XSTDFILL73_1816 VDD VSS sg13g2_FILL8
XSTDFILL73_1824 VDD VSS sg13g2_FILL8
XSTDFILL73_1832 VDD VSS sg13g2_FILL8
XSTDFILL73_1840 VDD VSS sg13g2_FILL8
XSTDFILL73_1848 VDD VSS sg13g2_FILL8
XSTDFILL73_1856 VDD VSS sg13g2_FILL8
XSTDFILL73_1864 VDD VSS sg13g2_FILL8
XSTDFILL73_1872 VDD VSS sg13g2_FILL8
XSTDFILL73_1880 VDD VSS sg13g2_FILL8
XSTDFILL73_1888 VDD VSS sg13g2_FILL8
XSTDFILL73_1896 VDD VSS sg13g2_FILL8
XSTDFILL73_1904 VDD VSS sg13g2_FILL8
XSTDFILL73_1912 VDD VSS sg13g2_FILL8
XSTDFILL73_1920 VDD VSS sg13g2_FILL8
XSTDFILL73_1928 VDD VSS sg13g2_FILL8
XSTDFILL73_1936 VDD VSS sg13g2_FILL8
XSTDFILL73_1944 VDD VSS sg13g2_FILL8
XSTDFILL73_1952 VDD VSS sg13g2_FILL8
XSTDFILL73_1960 VDD VSS sg13g2_FILL8
XSTDFILL73_1968 VDD VSS sg13g2_FILL8
XSTDFILL73_1976 VDD VSS sg13g2_FILL8
XSTDFILL73_1984 VDD VSS sg13g2_FILL8
XSTDFILL73_1992 VDD VSS sg13g2_FILL8
XSTDFILL73_2000 VDD VSS sg13g2_FILL8
XSTDFILL73_2008 VDD VSS sg13g2_FILL8
XSTDFILL73_2016 VDD VSS sg13g2_FILL8
XSTDFILL73_2024 VDD VSS sg13g2_FILL8
XSTDFILL73_2032 VDD VSS sg13g2_FILL8
XSTDFILL73_2040 VDD VSS sg13g2_FILL8
XSTDFILL73_2048 VDD VSS sg13g2_FILL8
XSTDFILL73_2056 VDD VSS sg13g2_FILL8
XSTDFILL73_2064 VDD VSS sg13g2_FILL8
XSTDFILL73_2072 VDD VSS sg13g2_FILL8
XSTDFILL73_2080 VDD VSS sg13g2_FILL8
XSTDFILL73_2088 VDD VSS sg13g2_FILL8
XSTDFILL73_2096 VDD VSS sg13g2_FILL8
XSTDFILL73_2104 VDD VSS sg13g2_FILL8
XSTDFILL73_2112 VDD VSS sg13g2_FILL8
XSTDFILL73_2120 VDD VSS sg13g2_FILL8
XSTDFILL73_2128 VDD VSS sg13g2_FILL8
XSTDFILL73_2136 VDD VSS sg13g2_FILL8
XSTDFILL73_2144 VDD VSS sg13g2_FILL8
XSTDFILL73_2152 VDD VSS sg13g2_FILL8
XSTDFILL73_2160 VDD VSS sg13g2_FILL8
XSTDFILL73_2168 VDD VSS sg13g2_FILL4
XSTDFILL74_0 VDD VSS sg13g2_FILL8
XSTDFILL74_8 VDD VSS sg13g2_FILL8
XSTDFILL74_16 VDD VSS sg13g2_FILL8
XSTDFILL74_24 VDD VSS sg13g2_FILL8
XSTDFILL74_32 VDD VSS sg13g2_FILL8
XSTDFILL74_40 VDD VSS sg13g2_FILL8
XSTDFILL74_48 VDD VSS sg13g2_FILL8
XSTDFILL74_56 VDD VSS sg13g2_FILL8
XSTDFILL74_64 VDD VSS sg13g2_FILL8
XSTDFILL74_72 VDD VSS sg13g2_FILL8
XSTDFILL74_80 VDD VSS sg13g2_FILL8
XSTDFILL74_88 VDD VSS sg13g2_FILL8
XSTDFILL74_96 VDD VSS sg13g2_FILL8
XSTDFILL74_104 VDD VSS sg13g2_FILL8
XSTDFILL74_112 VDD VSS sg13g2_FILL8
XSTDFILL74_120 VDD VSS sg13g2_FILL8
XSTDFILL74_128 VDD VSS sg13g2_FILL8
XSTDFILL74_136 VDD VSS sg13g2_FILL8
XSTDFILL74_144 VDD VSS sg13g2_FILL8
XSTDFILL74_152 VDD VSS sg13g2_FILL8
XSTDFILL74_160 VDD VSS sg13g2_FILL8
XSTDFILL74_168 VDD VSS sg13g2_FILL8
XSTDFILL74_176 VDD VSS sg13g2_FILL8
XSTDFILL74_184 VDD VSS sg13g2_FILL8
XSTDFILL74_192 VDD VSS sg13g2_FILL8
XSTDFILL74_200 VDD VSS sg13g2_FILL8
XSTDFILL74_208 VDD VSS sg13g2_FILL8
XSTDFILL74_216 VDD VSS sg13g2_FILL8
XSTDFILL74_224 VDD VSS sg13g2_FILL8
XSTDFILL74_232 VDD VSS sg13g2_FILL8
XSTDFILL74_240 VDD VSS sg13g2_FILL8
XSTDFILL74_248 VDD VSS sg13g2_FILL8
XSTDFILL74_256 VDD VSS sg13g2_FILL8
XSTDFILL74_264 VDD VSS sg13g2_FILL8
XSTDFILL74_272 VDD VSS sg13g2_FILL8
XSTDFILL74_280 VDD VSS sg13g2_FILL8
XSTDFILL74_288 VDD VSS sg13g2_FILL8
XSTDFILL74_296 VDD VSS sg13g2_FILL8
XSTDFILL74_304 VDD VSS sg13g2_FILL8
XSTDFILL74_312 VDD VSS sg13g2_FILL8
XSTDFILL74_320 VDD VSS sg13g2_FILL8
XSTDFILL74_328 VDD VSS sg13g2_FILL8
XSTDFILL74_336 VDD VSS sg13g2_FILL8
XSTDFILL74_344 VDD VSS sg13g2_FILL8
XSTDFILL74_352 VDD VSS sg13g2_FILL8
XSTDFILL74_360 VDD VSS sg13g2_FILL8
XSTDFILL74_368 VDD VSS sg13g2_FILL8
XSTDFILL74_376 VDD VSS sg13g2_FILL8
XSTDFILL74_384 VDD VSS sg13g2_FILL8
XSTDFILL74_392 VDD VSS sg13g2_FILL8
XSTDFILL74_400 VDD VSS sg13g2_FILL8
XSTDFILL74_408 VDD VSS sg13g2_FILL8
XSTDFILL74_416 VDD VSS sg13g2_FILL8
XSTDFILL74_424 VDD VSS sg13g2_FILL8
XSTDFILL74_432 VDD VSS sg13g2_FILL8
XSTDFILL74_440 VDD VSS sg13g2_FILL8
XSTDFILL74_448 VDD VSS sg13g2_FILL8
XSTDFILL74_456 VDD VSS sg13g2_FILL8
XSTDFILL74_464 VDD VSS sg13g2_FILL8
XSTDFILL74_472 VDD VSS sg13g2_FILL8
XSTDFILL74_480 VDD VSS sg13g2_FILL8
XSTDFILL74_488 VDD VSS sg13g2_FILL8
XSTDFILL74_496 VDD VSS sg13g2_FILL8
XSTDFILL74_504 VDD VSS sg13g2_FILL8
XSTDFILL74_512 VDD VSS sg13g2_FILL8
XSTDFILL74_520 VDD VSS sg13g2_FILL8
XSTDFILL74_528 VDD VSS sg13g2_FILL8
XSTDFILL74_536 VDD VSS sg13g2_FILL8
XSTDFILL74_544 VDD VSS sg13g2_FILL8
XSTDFILL74_552 VDD VSS sg13g2_FILL8
XSTDFILL74_560 VDD VSS sg13g2_FILL8
XSTDFILL74_568 VDD VSS sg13g2_FILL8
XSTDFILL74_576 VDD VSS sg13g2_FILL8
XSTDFILL74_584 VDD VSS sg13g2_FILL8
XSTDFILL74_592 VDD VSS sg13g2_FILL8
XSTDFILL74_600 VDD VSS sg13g2_FILL8
XSTDFILL74_608 VDD VSS sg13g2_FILL8
XSTDFILL74_616 VDD VSS sg13g2_FILL8
XSTDFILL74_624 VDD VSS sg13g2_FILL8
XSTDFILL74_632 VDD VSS sg13g2_FILL8
XSTDFILL74_640 VDD VSS sg13g2_FILL8
XSTDFILL74_648 VDD VSS sg13g2_FILL8
XSTDFILL74_656 VDD VSS sg13g2_FILL8
XSTDFILL74_664 VDD VSS sg13g2_FILL8
XSTDFILL74_672 VDD VSS sg13g2_FILL8
XSTDFILL74_680 VDD VSS sg13g2_FILL8
XSTDFILL74_688 VDD VSS sg13g2_FILL8
XSTDFILL74_696 VDD VSS sg13g2_FILL8
XSTDFILL74_704 VDD VSS sg13g2_FILL8
XSTDFILL74_712 VDD VSS sg13g2_FILL8
XSTDFILL74_720 VDD VSS sg13g2_FILL8
XSTDFILL74_728 VDD VSS sg13g2_FILL8
XSTDFILL74_736 VDD VSS sg13g2_FILL8
XSTDFILL74_744 VDD VSS sg13g2_FILL8
XSTDFILL74_752 VDD VSS sg13g2_FILL8
XSTDFILL74_760 VDD VSS sg13g2_FILL8
XSTDFILL74_768 VDD VSS sg13g2_FILL8
XSTDFILL74_776 VDD VSS sg13g2_FILL8
XSTDFILL74_784 VDD VSS sg13g2_FILL8
XSTDFILL74_792 VDD VSS sg13g2_FILL8
XSTDFILL74_800 VDD VSS sg13g2_FILL8
XSTDFILL74_808 VDD VSS sg13g2_FILL8
XSTDFILL74_816 VDD VSS sg13g2_FILL8
XSTDFILL74_824 VDD VSS sg13g2_FILL8
XSTDFILL74_832 VDD VSS sg13g2_FILL8
XSTDFILL74_840 VDD VSS sg13g2_FILL8
XSTDFILL74_848 VDD VSS sg13g2_FILL8
XSTDFILL74_856 VDD VSS sg13g2_FILL8
XSTDFILL74_864 VDD VSS sg13g2_FILL8
XSTDFILL74_872 VDD VSS sg13g2_FILL8
XSTDFILL74_880 VDD VSS sg13g2_FILL8
XSTDFILL74_888 VDD VSS sg13g2_FILL8
XSTDFILL74_896 VDD VSS sg13g2_FILL8
XSTDFILL74_904 VDD VSS sg13g2_FILL8
XSTDFILL74_912 VDD VSS sg13g2_FILL8
XSTDFILL74_920 VDD VSS sg13g2_FILL8
XSTDFILL74_928 VDD VSS sg13g2_FILL8
XSTDFILL74_936 VDD VSS sg13g2_FILL8
XSTDFILL74_944 VDD VSS sg13g2_FILL8
XSTDFILL74_952 VDD VSS sg13g2_FILL8
XSTDFILL74_960 VDD VSS sg13g2_FILL8
XSTDFILL74_968 VDD VSS sg13g2_FILL8
XSTDFILL74_976 VDD VSS sg13g2_FILL8
XSTDFILL74_984 VDD VSS sg13g2_FILL8
XSTDFILL74_992 VDD VSS sg13g2_FILL8
XSTDFILL74_1000 VDD VSS sg13g2_FILL8
XSTDFILL74_1008 VDD VSS sg13g2_FILL8
XSTDFILL74_1016 VDD VSS sg13g2_FILL8
XSTDFILL74_1024 VDD VSS sg13g2_FILL8
XSTDFILL74_1032 VDD VSS sg13g2_FILL8
XSTDFILL74_1040 VDD VSS sg13g2_FILL8
XSTDFILL74_1048 VDD VSS sg13g2_FILL8
XSTDFILL74_1056 VDD VSS sg13g2_FILL8
XSTDFILL74_1064 VDD VSS sg13g2_FILL8
XSTDFILL74_1072 VDD VSS sg13g2_FILL8
XSTDFILL74_1080 VDD VSS sg13g2_FILL8
XSTDFILL74_1088 VDD VSS sg13g2_FILL8
XSTDFILL74_1096 VDD VSS sg13g2_FILL8
XSTDFILL74_1104 VDD VSS sg13g2_FILL8
XSTDFILL74_1112 VDD VSS sg13g2_FILL8
XSTDFILL74_1120 VDD VSS sg13g2_FILL8
XSTDFILL74_1128 VDD VSS sg13g2_FILL8
XSTDFILL74_1136 VDD VSS sg13g2_FILL8
XSTDFILL74_1144 VDD VSS sg13g2_FILL8
XSTDFILL74_1152 VDD VSS sg13g2_FILL8
XSTDFILL74_1160 VDD VSS sg13g2_FILL8
XSTDFILL74_1168 VDD VSS sg13g2_FILL8
XSTDFILL74_1176 VDD VSS sg13g2_FILL8
XSTDFILL74_1184 VDD VSS sg13g2_FILL8
XSTDFILL74_1192 VDD VSS sg13g2_FILL8
XSTDFILL74_1200 VDD VSS sg13g2_FILL8
XSTDFILL74_1208 VDD VSS sg13g2_FILL8
XSTDFILL74_1216 VDD VSS sg13g2_FILL8
XSTDFILL74_1224 VDD VSS sg13g2_FILL8
XSTDFILL74_1232 VDD VSS sg13g2_FILL8
XSTDFILL74_1240 VDD VSS sg13g2_FILL8
XSTDFILL74_1248 VDD VSS sg13g2_FILL8
XSTDFILL74_1256 VDD VSS sg13g2_FILL8
XSTDFILL74_1264 VDD VSS sg13g2_FILL8
XSTDFILL74_1272 VDD VSS sg13g2_FILL8
XSTDFILL74_1280 VDD VSS sg13g2_FILL8
XSTDFILL74_1288 VDD VSS sg13g2_FILL8
XSTDFILL74_1296 VDD VSS sg13g2_FILL8
XSTDFILL74_1304 VDD VSS sg13g2_FILL8
XSTDFILL74_1312 VDD VSS sg13g2_FILL8
XSTDFILL74_1320 VDD VSS sg13g2_FILL8
XSTDFILL74_1328 VDD VSS sg13g2_FILL8
XSTDFILL74_1336 VDD VSS sg13g2_FILL8
XSTDFILL74_1344 VDD VSS sg13g2_FILL8
XSTDFILL74_1352 VDD VSS sg13g2_FILL8
XSTDFILL74_1360 VDD VSS sg13g2_FILL8
XSTDFILL74_1368 VDD VSS sg13g2_FILL8
XSTDFILL74_1376 VDD VSS sg13g2_FILL8
XSTDFILL74_1384 VDD VSS sg13g2_FILL8
XSTDFILL74_1392 VDD VSS sg13g2_FILL8
XSTDFILL74_1400 VDD VSS sg13g2_FILL8
XSTDFILL74_1408 VDD VSS sg13g2_FILL8
XSTDFILL74_1416 VDD VSS sg13g2_FILL8
XSTDFILL74_1424 VDD VSS sg13g2_FILL8
XSTDFILL74_1432 VDD VSS sg13g2_FILL8
XSTDFILL74_1440 VDD VSS sg13g2_FILL8
XSTDFILL74_1448 VDD VSS sg13g2_FILL8
XSTDFILL74_1456 VDD VSS sg13g2_FILL8
XSTDFILL74_1464 VDD VSS sg13g2_FILL8
XSTDFILL74_1472 VDD VSS sg13g2_FILL8
XSTDFILL74_1480 VDD VSS sg13g2_FILL8
XSTDFILL74_1488 VDD VSS sg13g2_FILL8
XSTDFILL74_1496 VDD VSS sg13g2_FILL8
XSTDFILL74_1504 VDD VSS sg13g2_FILL8
XSTDFILL74_1512 VDD VSS sg13g2_FILL8
XSTDFILL74_1520 VDD VSS sg13g2_FILL8
XSTDFILL74_1528 VDD VSS sg13g2_FILL8
XSTDFILL74_1536 VDD VSS sg13g2_FILL8
XSTDFILL74_1544 VDD VSS sg13g2_FILL8
XSTDFILL74_1552 VDD VSS sg13g2_FILL8
XSTDFILL74_1560 VDD VSS sg13g2_FILL8
XSTDFILL74_1568 VDD VSS sg13g2_FILL8
XSTDFILL74_1576 VDD VSS sg13g2_FILL8
XSTDFILL74_1584 VDD VSS sg13g2_FILL8
XSTDFILL74_1592 VDD VSS sg13g2_FILL8
XSTDFILL74_1600 VDD VSS sg13g2_FILL8
XSTDFILL74_1608 VDD VSS sg13g2_FILL8
XSTDFILL74_1616 VDD VSS sg13g2_FILL8
XSTDFILL74_1624 VDD VSS sg13g2_FILL8
XSTDFILL74_1632 VDD VSS sg13g2_FILL8
XSTDFILL74_1640 VDD VSS sg13g2_FILL8
XSTDFILL74_1648 VDD VSS sg13g2_FILL8
XSTDFILL74_1656 VDD VSS sg13g2_FILL8
XSTDFILL74_1664 VDD VSS sg13g2_FILL8
XSTDFILL74_1672 VDD VSS sg13g2_FILL8
XSTDFILL74_1680 VDD VSS sg13g2_FILL8
XSTDFILL74_1688 VDD VSS sg13g2_FILL8
XSTDFILL74_1696 VDD VSS sg13g2_FILL8
XSTDFILL74_1704 VDD VSS sg13g2_FILL8
XSTDFILL74_1712 VDD VSS sg13g2_FILL8
XSTDFILL74_1720 VDD VSS sg13g2_FILL8
XSTDFILL74_1728 VDD VSS sg13g2_FILL8
XSTDFILL74_1736 VDD VSS sg13g2_FILL8
XSTDFILL74_1744 VDD VSS sg13g2_FILL8
XSTDFILL74_1752 VDD VSS sg13g2_FILL8
XSTDFILL74_1760 VDD VSS sg13g2_FILL8
XSTDFILL74_1768 VDD VSS sg13g2_FILL8
XSTDFILL74_1776 VDD VSS sg13g2_FILL8
XSTDFILL74_1784 VDD VSS sg13g2_FILL8
XSTDFILL74_1792 VDD VSS sg13g2_FILL8
XSTDFILL74_1800 VDD VSS sg13g2_FILL8
XSTDFILL74_1808 VDD VSS sg13g2_FILL8
XSTDFILL74_1816 VDD VSS sg13g2_FILL8
XSTDFILL74_1824 VDD VSS sg13g2_FILL4
XSTDFILL74_1828 VDD VSS sg13g2_FILL2
XSTDFILL74_1835 VDD VSS sg13g2_FILL4
XSTDFILL74_1839 VDD VSS sg13g2_FILL1
XSTDFILL74_1848 VDD VSS sg13g2_FILL4
XSTDFILL74_1852 VDD VSS sg13g2_FILL1
XSTDFILL74_1858 VDD VSS sg13g2_FILL8
XSTDFILL74_1866 VDD VSS sg13g2_FILL8
XSTDFILL74_1882 VDD VSS sg13g2_FILL2
XSTDFILL74_1884 VDD VSS sg13g2_FILL1
XSTDFILL74_1890 VDD VSS sg13g2_FILL1
XSTDFILL74_1896 VDD VSS sg13g2_FILL8
XSTDFILL74_1904 VDD VSS sg13g2_FILL8
XSTDFILL74_1912 VDD VSS sg13g2_FILL8
XSTDFILL74_1920 VDD VSS sg13g2_FILL8
XSTDFILL74_1928 VDD VSS sg13g2_FILL8
XSTDFILL74_1936 VDD VSS sg13g2_FILL8
XSTDFILL74_1944 VDD VSS sg13g2_FILL8
XSTDFILL74_1952 VDD VSS sg13g2_FILL8
XSTDFILL74_1960 VDD VSS sg13g2_FILL8
XSTDFILL74_1968 VDD VSS sg13g2_FILL8
XSTDFILL74_1976 VDD VSS sg13g2_FILL8
XSTDFILL74_1984 VDD VSS sg13g2_FILL8
XSTDFILL74_1992 VDD VSS sg13g2_FILL8
XSTDFILL74_2000 VDD VSS sg13g2_FILL8
XSTDFILL74_2008 VDD VSS sg13g2_FILL8
XSTDFILL74_2016 VDD VSS sg13g2_FILL8
XSTDFILL74_2024 VDD VSS sg13g2_FILL8
XSTDFILL74_2032 VDD VSS sg13g2_FILL8
XSTDFILL74_2040 VDD VSS sg13g2_FILL8
XSTDFILL74_2048 VDD VSS sg13g2_FILL8
XSTDFILL74_2056 VDD VSS sg13g2_FILL8
XSTDFILL74_2064 VDD VSS sg13g2_FILL8
XSTDFILL74_2072 VDD VSS sg13g2_FILL8
XSTDFILL74_2080 VDD VSS sg13g2_FILL8
XSTDFILL74_2088 VDD VSS sg13g2_FILL8
XSTDFILL74_2096 VDD VSS sg13g2_FILL8
XSTDFILL74_2104 VDD VSS sg13g2_FILL8
XSTDFILL74_2112 VDD VSS sg13g2_FILL8
XSTDFILL74_2120 VDD VSS sg13g2_FILL8
XSTDFILL74_2128 VDD VSS sg13g2_FILL8
XSTDFILL74_2136 VDD VSS sg13g2_FILL8
XSTDFILL74_2144 VDD VSS sg13g2_FILL8
XSTDFILL74_2152 VDD VSS sg13g2_FILL8
XSTDFILL74_2160 VDD VSS sg13g2_FILL8
XSTDFILL74_2168 VDD VSS sg13g2_FILL4
XSTDFILL75_0 VDD VSS sg13g2_FILL8
XSTDFILL75_8 VDD VSS sg13g2_FILL8
XSTDFILL75_16 VDD VSS sg13g2_FILL8
XSTDFILL75_24 VDD VSS sg13g2_FILL8
XSTDFILL75_32 VDD VSS sg13g2_FILL8
XSTDFILL75_40 VDD VSS sg13g2_FILL8
XSTDFILL75_48 VDD VSS sg13g2_FILL8
XSTDFILL75_56 VDD VSS sg13g2_FILL8
XSTDFILL75_64 VDD VSS sg13g2_FILL8
XSTDFILL75_72 VDD VSS sg13g2_FILL8
XSTDFILL75_80 VDD VSS sg13g2_FILL8
XSTDFILL75_88 VDD VSS sg13g2_FILL8
XSTDFILL75_96 VDD VSS sg13g2_FILL8
XSTDFILL75_104 VDD VSS sg13g2_FILL8
XSTDFILL75_112 VDD VSS sg13g2_FILL8
XSTDFILL75_120 VDD VSS sg13g2_FILL8
XSTDFILL75_128 VDD VSS sg13g2_FILL8
XSTDFILL75_136 VDD VSS sg13g2_FILL8
XSTDFILL75_144 VDD VSS sg13g2_FILL8
XSTDFILL75_152 VDD VSS sg13g2_FILL8
XSTDFILL75_160 VDD VSS sg13g2_FILL8
XSTDFILL75_168 VDD VSS sg13g2_FILL8
XSTDFILL75_176 VDD VSS sg13g2_FILL8
XSTDFILL75_184 VDD VSS sg13g2_FILL8
XSTDFILL75_192 VDD VSS sg13g2_FILL8
XSTDFILL75_200 VDD VSS sg13g2_FILL8
XSTDFILL75_208 VDD VSS sg13g2_FILL8
XSTDFILL75_216 VDD VSS sg13g2_FILL8
XSTDFILL75_224 VDD VSS sg13g2_FILL8
XSTDFILL75_232 VDD VSS sg13g2_FILL8
XSTDFILL75_240 VDD VSS sg13g2_FILL8
XSTDFILL75_248 VDD VSS sg13g2_FILL8
XSTDFILL75_256 VDD VSS sg13g2_FILL8
XSTDFILL75_264 VDD VSS sg13g2_FILL8
XSTDFILL75_272 VDD VSS sg13g2_FILL8
XSTDFILL75_280 VDD VSS sg13g2_FILL8
XSTDFILL75_288 VDD VSS sg13g2_FILL8
XSTDFILL75_296 VDD VSS sg13g2_FILL8
XSTDFILL75_304 VDD VSS sg13g2_FILL8
XSTDFILL75_312 VDD VSS sg13g2_FILL8
XSTDFILL75_320 VDD VSS sg13g2_FILL8
XSTDFILL75_328 VDD VSS sg13g2_FILL8
XSTDFILL75_336 VDD VSS sg13g2_FILL8
XSTDFILL75_344 VDD VSS sg13g2_FILL8
XSTDFILL75_352 VDD VSS sg13g2_FILL8
XSTDFILL75_360 VDD VSS sg13g2_FILL8
XSTDFILL75_368 VDD VSS sg13g2_FILL8
XSTDFILL75_376 VDD VSS sg13g2_FILL8
XSTDFILL75_384 VDD VSS sg13g2_FILL8
XSTDFILL75_392 VDD VSS sg13g2_FILL8
XSTDFILL75_400 VDD VSS sg13g2_FILL8
XSTDFILL75_408 VDD VSS sg13g2_FILL8
XSTDFILL75_416 VDD VSS sg13g2_FILL8
XSTDFILL75_424 VDD VSS sg13g2_FILL8
XSTDFILL75_432 VDD VSS sg13g2_FILL8
XSTDFILL75_440 VDD VSS sg13g2_FILL8
XSTDFILL75_448 VDD VSS sg13g2_FILL8
XSTDFILL75_456 VDD VSS sg13g2_FILL8
XSTDFILL75_464 VDD VSS sg13g2_FILL8
XSTDFILL75_472 VDD VSS sg13g2_FILL8
XSTDFILL75_480 VDD VSS sg13g2_FILL8
XSTDFILL75_488 VDD VSS sg13g2_FILL8
XSTDFILL75_496 VDD VSS sg13g2_FILL8
XSTDFILL75_504 VDD VSS sg13g2_FILL8
XSTDFILL75_512 VDD VSS sg13g2_FILL8
XSTDFILL75_520 VDD VSS sg13g2_FILL8
XSTDFILL75_528 VDD VSS sg13g2_FILL8
XSTDFILL75_536 VDD VSS sg13g2_FILL8
XSTDFILL75_544 VDD VSS sg13g2_FILL8
XSTDFILL75_552 VDD VSS sg13g2_FILL8
XSTDFILL75_560 VDD VSS sg13g2_FILL8
XSTDFILL75_568 VDD VSS sg13g2_FILL8
XSTDFILL75_576 VDD VSS sg13g2_FILL8
XSTDFILL75_584 VDD VSS sg13g2_FILL8
XSTDFILL75_592 VDD VSS sg13g2_FILL8
XSTDFILL75_600 VDD VSS sg13g2_FILL8
XSTDFILL75_608 VDD VSS sg13g2_FILL8
XSTDFILL75_616 VDD VSS sg13g2_FILL8
XSTDFILL75_624 VDD VSS sg13g2_FILL8
XSTDFILL75_632 VDD VSS sg13g2_FILL8
XSTDFILL75_640 VDD VSS sg13g2_FILL8
XSTDFILL75_648 VDD VSS sg13g2_FILL8
XSTDFILL75_656 VDD VSS sg13g2_FILL8
XSTDFILL75_664 VDD VSS sg13g2_FILL8
XSTDFILL75_672 VDD VSS sg13g2_FILL8
XSTDFILL75_680 VDD VSS sg13g2_FILL8
XSTDFILL75_688 VDD VSS sg13g2_FILL8
XSTDFILL75_696 VDD VSS sg13g2_FILL8
XSTDFILL75_704 VDD VSS sg13g2_FILL8
XSTDFILL75_712 VDD VSS sg13g2_FILL8
XSTDFILL75_720 VDD VSS sg13g2_FILL8
XSTDFILL75_728 VDD VSS sg13g2_FILL8
XSTDFILL75_736 VDD VSS sg13g2_FILL8
XSTDFILL75_744 VDD VSS sg13g2_FILL8
XSTDFILL75_752 VDD VSS sg13g2_FILL8
XSTDFILL75_760 VDD VSS sg13g2_FILL8
XSTDFILL75_768 VDD VSS sg13g2_FILL8
XSTDFILL75_776 VDD VSS sg13g2_FILL8
XSTDFILL75_784 VDD VSS sg13g2_FILL8
XSTDFILL75_792 VDD VSS sg13g2_FILL8
XSTDFILL75_800 VDD VSS sg13g2_FILL8
XSTDFILL75_808 VDD VSS sg13g2_FILL8
XSTDFILL75_816 VDD VSS sg13g2_FILL8
XSTDFILL75_824 VDD VSS sg13g2_FILL8
XSTDFILL75_832 VDD VSS sg13g2_FILL8
XSTDFILL75_840 VDD VSS sg13g2_FILL8
XSTDFILL75_848 VDD VSS sg13g2_FILL8
XSTDFILL75_856 VDD VSS sg13g2_FILL8
XSTDFILL75_864 VDD VSS sg13g2_FILL8
XSTDFILL75_872 VDD VSS sg13g2_FILL8
XSTDFILL75_880 VDD VSS sg13g2_FILL8
XSTDFILL75_888 VDD VSS sg13g2_FILL8
XSTDFILL75_896 VDD VSS sg13g2_FILL8
XSTDFILL75_904 VDD VSS sg13g2_FILL8
XSTDFILL75_912 VDD VSS sg13g2_FILL8
XSTDFILL75_920 VDD VSS sg13g2_FILL8
XSTDFILL75_928 VDD VSS sg13g2_FILL8
XSTDFILL75_936 VDD VSS sg13g2_FILL8
XSTDFILL75_944 VDD VSS sg13g2_FILL8
XSTDFILL75_952 VDD VSS sg13g2_FILL8
XSTDFILL75_960 VDD VSS sg13g2_FILL8
XSTDFILL75_968 VDD VSS sg13g2_FILL8
XSTDFILL75_976 VDD VSS sg13g2_FILL8
XSTDFILL75_984 VDD VSS sg13g2_FILL8
XSTDFILL75_992 VDD VSS sg13g2_FILL8
XSTDFILL75_1000 VDD VSS sg13g2_FILL8
XSTDFILL75_1008 VDD VSS sg13g2_FILL8
XSTDFILL75_1016 VDD VSS sg13g2_FILL8
XSTDFILL75_1024 VDD VSS sg13g2_FILL8
XSTDFILL75_1032 VDD VSS sg13g2_FILL8
XSTDFILL75_1040 VDD VSS sg13g2_FILL8
XSTDFILL75_1048 VDD VSS sg13g2_FILL8
XSTDFILL75_1056 VDD VSS sg13g2_FILL8
XSTDFILL75_1064 VDD VSS sg13g2_FILL8
XSTDFILL75_1072 VDD VSS sg13g2_FILL8
XSTDFILL75_1080 VDD VSS sg13g2_FILL8
XSTDFILL75_1088 VDD VSS sg13g2_FILL8
XSTDFILL75_1096 VDD VSS sg13g2_FILL8
XSTDFILL75_1104 VDD VSS sg13g2_FILL8
XSTDFILL75_1112 VDD VSS sg13g2_FILL8
XSTDFILL75_1120 VDD VSS sg13g2_FILL8
XSTDFILL75_1128 VDD VSS sg13g2_FILL8
XSTDFILL75_1136 VDD VSS sg13g2_FILL8
XSTDFILL75_1144 VDD VSS sg13g2_FILL8
XSTDFILL75_1152 VDD VSS sg13g2_FILL8
XSTDFILL75_1160 VDD VSS sg13g2_FILL8
XSTDFILL75_1168 VDD VSS sg13g2_FILL8
XSTDFILL75_1176 VDD VSS sg13g2_FILL8
XSTDFILL75_1184 VDD VSS sg13g2_FILL8
XSTDFILL75_1192 VDD VSS sg13g2_FILL8
XSTDFILL75_1200 VDD VSS sg13g2_FILL8
XSTDFILL75_1208 VDD VSS sg13g2_FILL8
XSTDFILL75_1216 VDD VSS sg13g2_FILL8
XSTDFILL75_1224 VDD VSS sg13g2_FILL8
XSTDFILL75_1232 VDD VSS sg13g2_FILL8
XSTDFILL75_1240 VDD VSS sg13g2_FILL8
XSTDFILL75_1248 VDD VSS sg13g2_FILL8
XSTDFILL75_1256 VDD VSS sg13g2_FILL8
XSTDFILL75_1264 VDD VSS sg13g2_FILL8
XSTDFILL75_1272 VDD VSS sg13g2_FILL8
XSTDFILL75_1280 VDD VSS sg13g2_FILL8
XSTDFILL75_1288 VDD VSS sg13g2_FILL8
XSTDFILL75_1296 VDD VSS sg13g2_FILL8
XSTDFILL75_1304 VDD VSS sg13g2_FILL8
XSTDFILL75_1312 VDD VSS sg13g2_FILL8
XSTDFILL75_1320 VDD VSS sg13g2_FILL8
XSTDFILL75_1328 VDD VSS sg13g2_FILL8
XSTDFILL75_1336 VDD VSS sg13g2_FILL8
XSTDFILL75_1344 VDD VSS sg13g2_FILL8
XSTDFILL75_1352 VDD VSS sg13g2_FILL8
XSTDFILL75_1360 VDD VSS sg13g2_FILL8
XSTDFILL75_1368 VDD VSS sg13g2_FILL8
XSTDFILL75_1376 VDD VSS sg13g2_FILL8
XSTDFILL75_1384 VDD VSS sg13g2_FILL8
XSTDFILL75_1392 VDD VSS sg13g2_FILL8
XSTDFILL75_1400 VDD VSS sg13g2_FILL8
XSTDFILL75_1408 VDD VSS sg13g2_FILL8
XSTDFILL75_1416 VDD VSS sg13g2_FILL8
XSTDFILL75_1424 VDD VSS sg13g2_FILL8
XSTDFILL75_1432 VDD VSS sg13g2_FILL8
XSTDFILL75_1440 VDD VSS sg13g2_FILL8
XSTDFILL75_1448 VDD VSS sg13g2_FILL8
XSTDFILL75_1456 VDD VSS sg13g2_FILL8
XSTDFILL75_1464 VDD VSS sg13g2_FILL8
XSTDFILL75_1472 VDD VSS sg13g2_FILL8
XSTDFILL75_1480 VDD VSS sg13g2_FILL8
XSTDFILL75_1488 VDD VSS sg13g2_FILL8
XSTDFILL75_1496 VDD VSS sg13g2_FILL8
XSTDFILL75_1504 VDD VSS sg13g2_FILL8
XSTDFILL75_1512 VDD VSS sg13g2_FILL8
XSTDFILL75_1520 VDD VSS sg13g2_FILL8
XSTDFILL75_1528 VDD VSS sg13g2_FILL8
XSTDFILL75_1536 VDD VSS sg13g2_FILL8
XSTDFILL75_1544 VDD VSS sg13g2_FILL8
XSTDFILL75_1552 VDD VSS sg13g2_FILL8
XSTDFILL75_1560 VDD VSS sg13g2_FILL8
XSTDFILL75_1568 VDD VSS sg13g2_FILL8
XSTDFILL75_1576 VDD VSS sg13g2_FILL8
XSTDFILL75_1584 VDD VSS sg13g2_FILL8
XSTDFILL75_1592 VDD VSS sg13g2_FILL8
XSTDFILL75_1600 VDD VSS sg13g2_FILL8
XSTDFILL75_1608 VDD VSS sg13g2_FILL8
XSTDFILL75_1616 VDD VSS sg13g2_FILL8
XSTDFILL75_1624 VDD VSS sg13g2_FILL8
XSTDFILL75_1632 VDD VSS sg13g2_FILL8
XSTDFILL75_1640 VDD VSS sg13g2_FILL8
XSTDFILL75_1648 VDD VSS sg13g2_FILL8
XSTDFILL75_1656 VDD VSS sg13g2_FILL8
XSTDFILL75_1664 VDD VSS sg13g2_FILL8
XSTDFILL75_1672 VDD VSS sg13g2_FILL8
XSTDFILL75_1680 VDD VSS sg13g2_FILL8
XSTDFILL75_1688 VDD VSS sg13g2_FILL8
XSTDFILL75_1696 VDD VSS sg13g2_FILL8
XSTDFILL75_1704 VDD VSS sg13g2_FILL8
XSTDFILL75_1712 VDD VSS sg13g2_FILL8
XSTDFILL75_1720 VDD VSS sg13g2_FILL8
XSTDFILL75_1733 VDD VSS sg13g2_FILL8
XSTDFILL75_1741 VDD VSS sg13g2_FILL8
XSTDFILL75_1749 VDD VSS sg13g2_FILL2
XSTDFILL75_1772 VDD VSS sg13g2_FILL8
XSTDFILL75_1780 VDD VSS sg13g2_FILL1
XSTDFILL75_1807 VDD VSS sg13g2_FILL1
XSTDFILL75_1831 VDD VSS sg13g2_FILL2
XSTDFILL75_1846 VDD VSS sg13g2_FILL4
XSTDFILL75_1881 VDD VSS sg13g2_FILL2
XSTDFILL75_1883 VDD VSS sg13g2_FILL1
XSTDFILL75_1892 VDD VSS sg13g2_FILL4
XSTDFILL75_1941 VDD VSS sg13g2_FILL2
XSTDFILL75_1943 VDD VSS sg13g2_FILL1
XSTDFILL75_1967 VDD VSS sg13g2_FILL2
XSTDFILL75_1995 VDD VSS sg13g2_FILL2
XSTDFILL75_1997 VDD VSS sg13g2_FILL1
XSTDFILL75_2006 VDD VSS sg13g2_FILL8
XSTDFILL75_2014 VDD VSS sg13g2_FILL1
XSTDFILL75_2020 VDD VSS sg13g2_FILL1
XSTDFILL75_2034 VDD VSS sg13g2_FILL8
XSTDFILL75_2052 VDD VSS sg13g2_FILL8
XSTDFILL75_2060 VDD VSS sg13g2_FILL8
XSTDFILL75_2068 VDD VSS sg13g2_FILL8
XSTDFILL75_2076 VDD VSS sg13g2_FILL8
XSTDFILL75_2084 VDD VSS sg13g2_FILL8
XSTDFILL75_2092 VDD VSS sg13g2_FILL8
XSTDFILL75_2100 VDD VSS sg13g2_FILL8
XSTDFILL75_2108 VDD VSS sg13g2_FILL8
XSTDFILL75_2116 VDD VSS sg13g2_FILL8
XSTDFILL75_2124 VDD VSS sg13g2_FILL8
XSTDFILL75_2132 VDD VSS sg13g2_FILL8
XSTDFILL75_2140 VDD VSS sg13g2_FILL8
XSTDFILL75_2148 VDD VSS sg13g2_FILL8
XSTDFILL75_2156 VDD VSS sg13g2_FILL8
XSTDFILL75_2164 VDD VSS sg13g2_FILL8
XSTDFILL76_0 VDD VSS sg13g2_FILL8
XSTDFILL76_8 VDD VSS sg13g2_FILL8
XSTDFILL76_16 VDD VSS sg13g2_FILL8
XSTDFILL76_24 VDD VSS sg13g2_FILL8
XSTDFILL76_32 VDD VSS sg13g2_FILL8
XSTDFILL76_40 VDD VSS sg13g2_FILL8
XSTDFILL76_48 VDD VSS sg13g2_FILL8
XSTDFILL76_56 VDD VSS sg13g2_FILL8
XSTDFILL76_64 VDD VSS sg13g2_FILL8
XSTDFILL76_72 VDD VSS sg13g2_FILL8
XSTDFILL76_80 VDD VSS sg13g2_FILL8
XSTDFILL76_88 VDD VSS sg13g2_FILL8
XSTDFILL76_96 VDD VSS sg13g2_FILL8
XSTDFILL76_104 VDD VSS sg13g2_FILL8
XSTDFILL76_112 VDD VSS sg13g2_FILL8
XSTDFILL76_120 VDD VSS sg13g2_FILL8
XSTDFILL76_128 VDD VSS sg13g2_FILL8
XSTDFILL76_136 VDD VSS sg13g2_FILL8
XSTDFILL76_144 VDD VSS sg13g2_FILL8
XSTDFILL76_152 VDD VSS sg13g2_FILL8
XSTDFILL76_160 VDD VSS sg13g2_FILL8
XSTDFILL76_168 VDD VSS sg13g2_FILL8
XSTDFILL76_176 VDD VSS sg13g2_FILL8
XSTDFILL76_184 VDD VSS sg13g2_FILL8
XSTDFILL76_192 VDD VSS sg13g2_FILL8
XSTDFILL76_200 VDD VSS sg13g2_FILL8
XSTDFILL76_208 VDD VSS sg13g2_FILL8
XSTDFILL76_216 VDD VSS sg13g2_FILL8
XSTDFILL76_224 VDD VSS sg13g2_FILL8
XSTDFILL76_232 VDD VSS sg13g2_FILL8
XSTDFILL76_240 VDD VSS sg13g2_FILL8
XSTDFILL76_248 VDD VSS sg13g2_FILL8
XSTDFILL76_256 VDD VSS sg13g2_FILL8
XSTDFILL76_264 VDD VSS sg13g2_FILL8
XSTDFILL76_272 VDD VSS sg13g2_FILL8
XSTDFILL76_280 VDD VSS sg13g2_FILL8
XSTDFILL76_288 VDD VSS sg13g2_FILL8
XSTDFILL76_296 VDD VSS sg13g2_FILL8
XSTDFILL76_304 VDD VSS sg13g2_FILL8
XSTDFILL76_312 VDD VSS sg13g2_FILL8
XSTDFILL76_320 VDD VSS sg13g2_FILL8
XSTDFILL76_328 VDD VSS sg13g2_FILL8
XSTDFILL76_336 VDD VSS sg13g2_FILL8
XSTDFILL76_344 VDD VSS sg13g2_FILL8
XSTDFILL76_352 VDD VSS sg13g2_FILL8
XSTDFILL76_360 VDD VSS sg13g2_FILL8
XSTDFILL76_368 VDD VSS sg13g2_FILL8
XSTDFILL76_376 VDD VSS sg13g2_FILL8
XSTDFILL76_384 VDD VSS sg13g2_FILL8
XSTDFILL76_392 VDD VSS sg13g2_FILL8
XSTDFILL76_400 VDD VSS sg13g2_FILL8
XSTDFILL76_408 VDD VSS sg13g2_FILL8
XSTDFILL76_416 VDD VSS sg13g2_FILL8
XSTDFILL76_424 VDD VSS sg13g2_FILL8
XSTDFILL76_432 VDD VSS sg13g2_FILL8
XSTDFILL76_440 VDD VSS sg13g2_FILL8
XSTDFILL76_448 VDD VSS sg13g2_FILL8
XSTDFILL76_456 VDD VSS sg13g2_FILL8
XSTDFILL76_464 VDD VSS sg13g2_FILL8
XSTDFILL76_472 VDD VSS sg13g2_FILL8
XSTDFILL76_480 VDD VSS sg13g2_FILL8
XSTDFILL76_488 VDD VSS sg13g2_FILL8
XSTDFILL76_496 VDD VSS sg13g2_FILL8
XSTDFILL76_504 VDD VSS sg13g2_FILL8
XSTDFILL76_512 VDD VSS sg13g2_FILL8
XSTDFILL76_520 VDD VSS sg13g2_FILL8
XSTDFILL76_528 VDD VSS sg13g2_FILL8
XSTDFILL76_536 VDD VSS sg13g2_FILL8
XSTDFILL76_544 VDD VSS sg13g2_FILL8
XSTDFILL76_552 VDD VSS sg13g2_FILL8
XSTDFILL76_560 VDD VSS sg13g2_FILL8
XSTDFILL76_568 VDD VSS sg13g2_FILL8
XSTDFILL76_576 VDD VSS sg13g2_FILL8
XSTDFILL76_584 VDD VSS sg13g2_FILL8
XSTDFILL76_592 VDD VSS sg13g2_FILL8
XSTDFILL76_600 VDD VSS sg13g2_FILL8
XSTDFILL76_608 VDD VSS sg13g2_FILL8
XSTDFILL76_616 VDD VSS sg13g2_FILL8
XSTDFILL76_624 VDD VSS sg13g2_FILL8
XSTDFILL76_632 VDD VSS sg13g2_FILL8
XSTDFILL76_640 VDD VSS sg13g2_FILL8
XSTDFILL76_648 VDD VSS sg13g2_FILL8
XSTDFILL76_656 VDD VSS sg13g2_FILL8
XSTDFILL76_664 VDD VSS sg13g2_FILL8
XSTDFILL76_672 VDD VSS sg13g2_FILL8
XSTDFILL76_680 VDD VSS sg13g2_FILL8
XSTDFILL76_688 VDD VSS sg13g2_FILL8
XSTDFILL76_696 VDD VSS sg13g2_FILL8
XSTDFILL76_704 VDD VSS sg13g2_FILL8
XSTDFILL76_712 VDD VSS sg13g2_FILL8
XSTDFILL76_720 VDD VSS sg13g2_FILL8
XSTDFILL76_728 VDD VSS sg13g2_FILL8
XSTDFILL76_736 VDD VSS sg13g2_FILL8
XSTDFILL76_744 VDD VSS sg13g2_FILL8
XSTDFILL76_752 VDD VSS sg13g2_FILL8
XSTDFILL76_760 VDD VSS sg13g2_FILL8
XSTDFILL76_768 VDD VSS sg13g2_FILL8
XSTDFILL76_776 VDD VSS sg13g2_FILL8
XSTDFILL76_784 VDD VSS sg13g2_FILL8
XSTDFILL76_792 VDD VSS sg13g2_FILL8
XSTDFILL76_800 VDD VSS sg13g2_FILL8
XSTDFILL76_808 VDD VSS sg13g2_FILL8
XSTDFILL76_816 VDD VSS sg13g2_FILL8
XSTDFILL76_824 VDD VSS sg13g2_FILL8
XSTDFILL76_832 VDD VSS sg13g2_FILL8
XSTDFILL76_840 VDD VSS sg13g2_FILL8
XSTDFILL76_848 VDD VSS sg13g2_FILL8
XSTDFILL76_856 VDD VSS sg13g2_FILL8
XSTDFILL76_864 VDD VSS sg13g2_FILL8
XSTDFILL76_872 VDD VSS sg13g2_FILL8
XSTDFILL76_880 VDD VSS sg13g2_FILL8
XSTDFILL76_888 VDD VSS sg13g2_FILL8
XSTDFILL76_896 VDD VSS sg13g2_FILL8
XSTDFILL76_904 VDD VSS sg13g2_FILL8
XSTDFILL76_912 VDD VSS sg13g2_FILL8
XSTDFILL76_920 VDD VSS sg13g2_FILL8
XSTDFILL76_928 VDD VSS sg13g2_FILL8
XSTDFILL76_936 VDD VSS sg13g2_FILL8
XSTDFILL76_944 VDD VSS sg13g2_FILL8
XSTDFILL76_952 VDD VSS sg13g2_FILL8
XSTDFILL76_960 VDD VSS sg13g2_FILL8
XSTDFILL76_968 VDD VSS sg13g2_FILL8
XSTDFILL76_976 VDD VSS sg13g2_FILL8
XSTDFILL76_984 VDD VSS sg13g2_FILL8
XSTDFILL76_992 VDD VSS sg13g2_FILL8
XSTDFILL76_1000 VDD VSS sg13g2_FILL8
XSTDFILL76_1008 VDD VSS sg13g2_FILL8
XSTDFILL76_1016 VDD VSS sg13g2_FILL8
XSTDFILL76_1024 VDD VSS sg13g2_FILL8
XSTDFILL76_1032 VDD VSS sg13g2_FILL8
XSTDFILL76_1040 VDD VSS sg13g2_FILL8
XSTDFILL76_1048 VDD VSS sg13g2_FILL8
XSTDFILL76_1056 VDD VSS sg13g2_FILL8
XSTDFILL76_1064 VDD VSS sg13g2_FILL8
XSTDFILL76_1072 VDD VSS sg13g2_FILL8
XSTDFILL76_1080 VDD VSS sg13g2_FILL8
XSTDFILL76_1088 VDD VSS sg13g2_FILL8
XSTDFILL76_1096 VDD VSS sg13g2_FILL8
XSTDFILL76_1104 VDD VSS sg13g2_FILL8
XSTDFILL76_1112 VDD VSS sg13g2_FILL8
XSTDFILL76_1120 VDD VSS sg13g2_FILL8
XSTDFILL76_1128 VDD VSS sg13g2_FILL8
XSTDFILL76_1136 VDD VSS sg13g2_FILL8
XSTDFILL76_1144 VDD VSS sg13g2_FILL8
XSTDFILL76_1152 VDD VSS sg13g2_FILL8
XSTDFILL76_1160 VDD VSS sg13g2_FILL8
XSTDFILL76_1168 VDD VSS sg13g2_FILL8
XSTDFILL76_1176 VDD VSS sg13g2_FILL8
XSTDFILL76_1184 VDD VSS sg13g2_FILL8
XSTDFILL76_1192 VDD VSS sg13g2_FILL8
XSTDFILL76_1200 VDD VSS sg13g2_FILL8
XSTDFILL76_1208 VDD VSS sg13g2_FILL8
XSTDFILL76_1216 VDD VSS sg13g2_FILL8
XSTDFILL76_1224 VDD VSS sg13g2_FILL8
XSTDFILL76_1232 VDD VSS sg13g2_FILL8
XSTDFILL76_1240 VDD VSS sg13g2_FILL8
XSTDFILL76_1248 VDD VSS sg13g2_FILL8
XSTDFILL76_1256 VDD VSS sg13g2_FILL8
XSTDFILL76_1264 VDD VSS sg13g2_FILL8
XSTDFILL76_1272 VDD VSS sg13g2_FILL8
XSTDFILL76_1280 VDD VSS sg13g2_FILL8
XSTDFILL76_1288 VDD VSS sg13g2_FILL8
XSTDFILL76_1296 VDD VSS sg13g2_FILL8
XSTDFILL76_1304 VDD VSS sg13g2_FILL8
XSTDFILL76_1312 VDD VSS sg13g2_FILL8
XSTDFILL76_1320 VDD VSS sg13g2_FILL8
XSTDFILL76_1328 VDD VSS sg13g2_FILL8
XSTDFILL76_1336 VDD VSS sg13g2_FILL8
XSTDFILL76_1344 VDD VSS sg13g2_FILL8
XSTDFILL76_1352 VDD VSS sg13g2_FILL8
XSTDFILL76_1360 VDD VSS sg13g2_FILL8
XSTDFILL76_1368 VDD VSS sg13g2_FILL8
XSTDFILL76_1376 VDD VSS sg13g2_FILL8
XSTDFILL76_1384 VDD VSS sg13g2_FILL8
XSTDFILL76_1392 VDD VSS sg13g2_FILL8
XSTDFILL76_1400 VDD VSS sg13g2_FILL8
XSTDFILL76_1408 VDD VSS sg13g2_FILL8
XSTDFILL76_1416 VDD VSS sg13g2_FILL8
XSTDFILL76_1424 VDD VSS sg13g2_FILL8
XSTDFILL76_1432 VDD VSS sg13g2_FILL8
XSTDFILL76_1440 VDD VSS sg13g2_FILL8
XSTDFILL76_1448 VDD VSS sg13g2_FILL8
XSTDFILL76_1456 VDD VSS sg13g2_FILL8
XSTDFILL76_1464 VDD VSS sg13g2_FILL8
XSTDFILL76_1472 VDD VSS sg13g2_FILL8
XSTDFILL76_1480 VDD VSS sg13g2_FILL8
XSTDFILL76_1488 VDD VSS sg13g2_FILL8
XSTDFILL76_1496 VDD VSS sg13g2_FILL8
XSTDFILL76_1504 VDD VSS sg13g2_FILL8
XSTDFILL76_1512 VDD VSS sg13g2_FILL8
XSTDFILL76_1520 VDD VSS sg13g2_FILL8
XSTDFILL76_1528 VDD VSS sg13g2_FILL2
XSTDFILL76_1530 VDD VSS sg13g2_FILL1
XSTDFILL77_0 VDD VSS sg13g2_FILL8
XSTDFILL77_8 VDD VSS sg13g2_FILL8
XSTDFILL77_16 VDD VSS sg13g2_FILL8
XSTDFILL77_24 VDD VSS sg13g2_FILL8
XSTDFILL77_32 VDD VSS sg13g2_FILL8
XSTDFILL77_40 VDD VSS sg13g2_FILL8
XSTDFILL77_48 VDD VSS sg13g2_FILL8
XSTDFILL77_56 VDD VSS sg13g2_FILL8
XSTDFILL77_64 VDD VSS sg13g2_FILL8
XSTDFILL77_72 VDD VSS sg13g2_FILL8
XSTDFILL77_80 VDD VSS sg13g2_FILL8
XSTDFILL77_88 VDD VSS sg13g2_FILL8
XSTDFILL77_96 VDD VSS sg13g2_FILL8
XSTDFILL77_104 VDD VSS sg13g2_FILL8
XSTDFILL77_112 VDD VSS sg13g2_FILL8
XSTDFILL77_120 VDD VSS sg13g2_FILL8
XSTDFILL77_128 VDD VSS sg13g2_FILL8
XSTDFILL77_136 VDD VSS sg13g2_FILL8
XSTDFILL77_144 VDD VSS sg13g2_FILL8
XSTDFILL77_152 VDD VSS sg13g2_FILL8
XSTDFILL77_160 VDD VSS sg13g2_FILL8
XSTDFILL77_168 VDD VSS sg13g2_FILL8
XSTDFILL77_176 VDD VSS sg13g2_FILL8
XSTDFILL77_184 VDD VSS sg13g2_FILL8
XSTDFILL77_192 VDD VSS sg13g2_FILL8
XSTDFILL77_200 VDD VSS sg13g2_FILL8
XSTDFILL77_208 VDD VSS sg13g2_FILL8
XSTDFILL77_216 VDD VSS sg13g2_FILL8
XSTDFILL77_224 VDD VSS sg13g2_FILL8
XSTDFILL77_232 VDD VSS sg13g2_FILL8
XSTDFILL77_240 VDD VSS sg13g2_FILL8
XSTDFILL77_248 VDD VSS sg13g2_FILL8
XSTDFILL77_256 VDD VSS sg13g2_FILL8
XSTDFILL77_264 VDD VSS sg13g2_FILL8
XSTDFILL77_272 VDD VSS sg13g2_FILL8
XSTDFILL77_280 VDD VSS sg13g2_FILL8
XSTDFILL77_288 VDD VSS sg13g2_FILL8
XSTDFILL77_296 VDD VSS sg13g2_FILL8
XSTDFILL77_304 VDD VSS sg13g2_FILL8
XSTDFILL77_312 VDD VSS sg13g2_FILL8
XSTDFILL77_320 VDD VSS sg13g2_FILL8
XSTDFILL77_328 VDD VSS sg13g2_FILL8
XSTDFILL77_336 VDD VSS sg13g2_FILL8
XSTDFILL77_344 VDD VSS sg13g2_FILL8
XSTDFILL77_352 VDD VSS sg13g2_FILL8
XSTDFILL77_360 VDD VSS sg13g2_FILL8
XSTDFILL77_368 VDD VSS sg13g2_FILL8
XSTDFILL77_376 VDD VSS sg13g2_FILL8
XSTDFILL77_384 VDD VSS sg13g2_FILL8
XSTDFILL77_392 VDD VSS sg13g2_FILL8
XSTDFILL77_400 VDD VSS sg13g2_FILL8
XSTDFILL77_408 VDD VSS sg13g2_FILL8
XSTDFILL77_416 VDD VSS sg13g2_FILL8
XSTDFILL77_424 VDD VSS sg13g2_FILL8
XSTDFILL77_432 VDD VSS sg13g2_FILL8
XSTDFILL77_440 VDD VSS sg13g2_FILL8
XSTDFILL77_448 VDD VSS sg13g2_FILL8
XSTDFILL77_456 VDD VSS sg13g2_FILL8
XSTDFILL77_464 VDD VSS sg13g2_FILL8
XSTDFILL77_472 VDD VSS sg13g2_FILL8
XSTDFILL77_480 VDD VSS sg13g2_FILL8
XSTDFILL77_488 VDD VSS sg13g2_FILL8
XSTDFILL77_496 VDD VSS sg13g2_FILL8
XSTDFILL77_504 VDD VSS sg13g2_FILL8
XSTDFILL77_512 VDD VSS sg13g2_FILL8
XSTDFILL77_520 VDD VSS sg13g2_FILL8
XSTDFILL77_528 VDD VSS sg13g2_FILL8
XSTDFILL77_536 VDD VSS sg13g2_FILL8
XSTDFILL77_544 VDD VSS sg13g2_FILL8
XSTDFILL77_552 VDD VSS sg13g2_FILL8
XSTDFILL77_560 VDD VSS sg13g2_FILL8
XSTDFILL77_568 VDD VSS sg13g2_FILL8
XSTDFILL77_576 VDD VSS sg13g2_FILL8
XSTDFILL77_584 VDD VSS sg13g2_FILL8
XSTDFILL77_592 VDD VSS sg13g2_FILL8
XSTDFILL77_600 VDD VSS sg13g2_FILL8
XSTDFILL77_608 VDD VSS sg13g2_FILL8
XSTDFILL77_616 VDD VSS sg13g2_FILL8
XSTDFILL77_624 VDD VSS sg13g2_FILL8
XSTDFILL77_632 VDD VSS sg13g2_FILL8
XSTDFILL77_640 VDD VSS sg13g2_FILL8
XSTDFILL77_648 VDD VSS sg13g2_FILL8
XSTDFILL77_656 VDD VSS sg13g2_FILL8
XSTDFILL77_664 VDD VSS sg13g2_FILL8
XSTDFILL77_672 VDD VSS sg13g2_FILL8
XSTDFILL77_680 VDD VSS sg13g2_FILL8
XSTDFILL77_688 VDD VSS sg13g2_FILL8
XSTDFILL77_696 VDD VSS sg13g2_FILL8
XSTDFILL77_704 VDD VSS sg13g2_FILL8
XSTDFILL77_712 VDD VSS sg13g2_FILL8
XSTDFILL77_720 VDD VSS sg13g2_FILL8
XSTDFILL77_728 VDD VSS sg13g2_FILL8
XSTDFILL77_736 VDD VSS sg13g2_FILL8
XSTDFILL77_744 VDD VSS sg13g2_FILL8
XSTDFILL77_752 VDD VSS sg13g2_FILL8
XSTDFILL77_760 VDD VSS sg13g2_FILL8
XSTDFILL77_768 VDD VSS sg13g2_FILL8
XSTDFILL77_776 VDD VSS sg13g2_FILL8
XSTDFILL77_784 VDD VSS sg13g2_FILL8
XSTDFILL77_792 VDD VSS sg13g2_FILL8
XSTDFILL77_800 VDD VSS sg13g2_FILL8
XSTDFILL77_808 VDD VSS sg13g2_FILL8
XSTDFILL77_816 VDD VSS sg13g2_FILL8
XSTDFILL77_824 VDD VSS sg13g2_FILL8
XSTDFILL77_832 VDD VSS sg13g2_FILL8
XSTDFILL77_840 VDD VSS sg13g2_FILL8
XSTDFILL77_848 VDD VSS sg13g2_FILL8
XSTDFILL77_856 VDD VSS sg13g2_FILL8
XSTDFILL77_864 VDD VSS sg13g2_FILL8
XSTDFILL77_872 VDD VSS sg13g2_FILL8
XSTDFILL77_880 VDD VSS sg13g2_FILL8
XSTDFILL77_888 VDD VSS sg13g2_FILL8
XSTDFILL77_896 VDD VSS sg13g2_FILL8
XSTDFILL77_904 VDD VSS sg13g2_FILL8
XSTDFILL77_912 VDD VSS sg13g2_FILL8
XSTDFILL77_920 VDD VSS sg13g2_FILL8
XSTDFILL77_928 VDD VSS sg13g2_FILL8
XSTDFILL77_936 VDD VSS sg13g2_FILL8
XSTDFILL77_944 VDD VSS sg13g2_FILL8
XSTDFILL77_952 VDD VSS sg13g2_FILL8
XSTDFILL77_960 VDD VSS sg13g2_FILL8
XSTDFILL77_968 VDD VSS sg13g2_FILL8
XSTDFILL77_976 VDD VSS sg13g2_FILL8
XSTDFILL77_984 VDD VSS sg13g2_FILL8
XSTDFILL77_992 VDD VSS sg13g2_FILL8
XSTDFILL77_1000 VDD VSS sg13g2_FILL8
XSTDFILL77_1008 VDD VSS sg13g2_FILL8
XSTDFILL77_1016 VDD VSS sg13g2_FILL8
XSTDFILL77_1024 VDD VSS sg13g2_FILL8
XSTDFILL77_1032 VDD VSS sg13g2_FILL8
XSTDFILL77_1040 VDD VSS sg13g2_FILL8
XSTDFILL77_1048 VDD VSS sg13g2_FILL8
XSTDFILL77_1056 VDD VSS sg13g2_FILL8
XSTDFILL77_1064 VDD VSS sg13g2_FILL8
XSTDFILL77_1072 VDD VSS sg13g2_FILL8
XSTDFILL77_1080 VDD VSS sg13g2_FILL8
XSTDFILL77_1088 VDD VSS sg13g2_FILL8
XSTDFILL77_1096 VDD VSS sg13g2_FILL8
XSTDFILL77_1104 VDD VSS sg13g2_FILL8
XSTDFILL77_1112 VDD VSS sg13g2_FILL8
XSTDFILL77_1120 VDD VSS sg13g2_FILL8
XSTDFILL77_1128 VDD VSS sg13g2_FILL8
XSTDFILL77_1136 VDD VSS sg13g2_FILL8
XSTDFILL77_1144 VDD VSS sg13g2_FILL8
XSTDFILL77_1152 VDD VSS sg13g2_FILL8
XSTDFILL77_1160 VDD VSS sg13g2_FILL8
XSTDFILL77_1168 VDD VSS sg13g2_FILL8
XSTDFILL77_1176 VDD VSS sg13g2_FILL8
XSTDFILL77_1184 VDD VSS sg13g2_FILL8
XSTDFILL77_1192 VDD VSS sg13g2_FILL8
XSTDFILL77_1200 VDD VSS sg13g2_FILL8
XSTDFILL77_1208 VDD VSS sg13g2_FILL8
XSTDFILL77_1216 VDD VSS sg13g2_FILL8
XSTDFILL77_1224 VDD VSS sg13g2_FILL8
XSTDFILL77_1232 VDD VSS sg13g2_FILL8
XSTDFILL77_1240 VDD VSS sg13g2_FILL8
XSTDFILL77_1248 VDD VSS sg13g2_FILL8
XSTDFILL77_1256 VDD VSS sg13g2_FILL8
XSTDFILL77_1264 VDD VSS sg13g2_FILL8
XSTDFILL77_1272 VDD VSS sg13g2_FILL8
XSTDFILL77_1280 VDD VSS sg13g2_FILL8
XSTDFILL77_1288 VDD VSS sg13g2_FILL8
XSTDFILL77_1296 VDD VSS sg13g2_FILL8
XSTDFILL77_1304 VDD VSS sg13g2_FILL8
XSTDFILL77_1312 VDD VSS sg13g2_FILL8
XSTDFILL77_1320 VDD VSS sg13g2_FILL8
XSTDFILL77_1328 VDD VSS sg13g2_FILL8
XSTDFILL77_1336 VDD VSS sg13g2_FILL8
XSTDFILL77_1344 VDD VSS sg13g2_FILL8
XSTDFILL77_1352 VDD VSS sg13g2_FILL8
XSTDFILL77_1360 VDD VSS sg13g2_FILL8
XSTDFILL77_1368 VDD VSS sg13g2_FILL8
XSTDFILL77_1376 VDD VSS sg13g2_FILL8
XSTDFILL77_1384 VDD VSS sg13g2_FILL8
XSTDFILL77_1392 VDD VSS sg13g2_FILL8
XSTDFILL77_1400 VDD VSS sg13g2_FILL8
XSTDFILL77_1408 VDD VSS sg13g2_FILL8
XSTDFILL77_1416 VDD VSS sg13g2_FILL8
XSTDFILL77_1424 VDD VSS sg13g2_FILL8
XSTDFILL77_1432 VDD VSS sg13g2_FILL8
XSTDFILL77_1440 VDD VSS sg13g2_FILL8
XSTDFILL77_1448 VDD VSS sg13g2_FILL8
XSTDFILL77_1456 VDD VSS sg13g2_FILL8
XSTDFILL77_1464 VDD VSS sg13g2_FILL8
XSTDFILL77_1472 VDD VSS sg13g2_FILL8
XSTDFILL77_1480 VDD VSS sg13g2_FILL8
XSTDFILL77_1488 VDD VSS sg13g2_FILL8
XSTDFILL77_1496 VDD VSS sg13g2_FILL8
XSTDFILL77_1504 VDD VSS sg13g2_FILL8
XSTDFILL77_1512 VDD VSS sg13g2_FILL8
XSTDFILL77_1520 VDD VSS sg13g2_FILL8
XSTDFILL77_1528 VDD VSS sg13g2_FILL2
XSTDFILL77_1530 VDD VSS sg13g2_FILL1
XSTDFILL78_0 VDD VSS sg13g2_FILL8
XSTDFILL78_8 VDD VSS sg13g2_FILL8
XSTDFILL78_16 VDD VSS sg13g2_FILL8
XSTDFILL78_24 VDD VSS sg13g2_FILL8
XSTDFILL78_32 VDD VSS sg13g2_FILL8
XSTDFILL78_40 VDD VSS sg13g2_FILL8
XSTDFILL78_48 VDD VSS sg13g2_FILL8
XSTDFILL78_56 VDD VSS sg13g2_FILL8
XSTDFILL78_64 VDD VSS sg13g2_FILL8
XSTDFILL78_72 VDD VSS sg13g2_FILL8
XSTDFILL78_80 VDD VSS sg13g2_FILL8
XSTDFILL78_88 VDD VSS sg13g2_FILL8
XSTDFILL78_96 VDD VSS sg13g2_FILL8
XSTDFILL78_104 VDD VSS sg13g2_FILL8
XSTDFILL78_112 VDD VSS sg13g2_FILL8
XSTDFILL78_120 VDD VSS sg13g2_FILL8
XSTDFILL78_128 VDD VSS sg13g2_FILL8
XSTDFILL78_136 VDD VSS sg13g2_FILL8
XSTDFILL78_144 VDD VSS sg13g2_FILL8
XSTDFILL78_152 VDD VSS sg13g2_FILL8
XSTDFILL78_160 VDD VSS sg13g2_FILL8
XSTDFILL78_168 VDD VSS sg13g2_FILL8
XSTDFILL78_176 VDD VSS sg13g2_FILL8
XSTDFILL78_184 VDD VSS sg13g2_FILL8
XSTDFILL78_192 VDD VSS sg13g2_FILL8
XSTDFILL78_200 VDD VSS sg13g2_FILL8
XSTDFILL78_208 VDD VSS sg13g2_FILL8
XSTDFILL78_216 VDD VSS sg13g2_FILL8
XSTDFILL78_224 VDD VSS sg13g2_FILL8
XSTDFILL78_232 VDD VSS sg13g2_FILL8
XSTDFILL78_240 VDD VSS sg13g2_FILL8
XSTDFILL78_248 VDD VSS sg13g2_FILL8
XSTDFILL78_256 VDD VSS sg13g2_FILL8
XSTDFILL78_264 VDD VSS sg13g2_FILL8
XSTDFILL78_272 VDD VSS sg13g2_FILL8
XSTDFILL78_280 VDD VSS sg13g2_FILL8
XSTDFILL78_288 VDD VSS sg13g2_FILL8
XSTDFILL78_296 VDD VSS sg13g2_FILL8
XSTDFILL78_304 VDD VSS sg13g2_FILL8
XSTDFILL78_312 VDD VSS sg13g2_FILL8
XSTDFILL78_320 VDD VSS sg13g2_FILL8
XSTDFILL78_328 VDD VSS sg13g2_FILL8
XSTDFILL78_336 VDD VSS sg13g2_FILL8
XSTDFILL78_344 VDD VSS sg13g2_FILL8
XSTDFILL78_352 VDD VSS sg13g2_FILL8
XSTDFILL78_360 VDD VSS sg13g2_FILL8
XSTDFILL78_368 VDD VSS sg13g2_FILL8
XSTDFILL78_376 VDD VSS sg13g2_FILL8
XSTDFILL78_384 VDD VSS sg13g2_FILL8
XSTDFILL78_392 VDD VSS sg13g2_FILL8
XSTDFILL78_400 VDD VSS sg13g2_FILL8
XSTDFILL78_408 VDD VSS sg13g2_FILL8
XSTDFILL78_416 VDD VSS sg13g2_FILL8
XSTDFILL78_424 VDD VSS sg13g2_FILL8
XSTDFILL78_432 VDD VSS sg13g2_FILL8
XSTDFILL78_440 VDD VSS sg13g2_FILL8
XSTDFILL78_448 VDD VSS sg13g2_FILL8
XSTDFILL78_456 VDD VSS sg13g2_FILL8
XSTDFILL78_464 VDD VSS sg13g2_FILL8
XSTDFILL78_472 VDD VSS sg13g2_FILL8
XSTDFILL78_480 VDD VSS sg13g2_FILL8
XSTDFILL78_488 VDD VSS sg13g2_FILL8
XSTDFILL78_496 VDD VSS sg13g2_FILL8
XSTDFILL78_504 VDD VSS sg13g2_FILL8
XSTDFILL78_512 VDD VSS sg13g2_FILL8
XSTDFILL78_520 VDD VSS sg13g2_FILL8
XSTDFILL78_528 VDD VSS sg13g2_FILL8
XSTDFILL78_536 VDD VSS sg13g2_FILL8
XSTDFILL78_544 VDD VSS sg13g2_FILL8
XSTDFILL78_552 VDD VSS sg13g2_FILL8
XSTDFILL78_560 VDD VSS sg13g2_FILL8
XSTDFILL78_568 VDD VSS sg13g2_FILL8
XSTDFILL78_576 VDD VSS sg13g2_FILL8
XSTDFILL78_584 VDD VSS sg13g2_FILL8
XSTDFILL78_592 VDD VSS sg13g2_FILL8
XSTDFILL78_600 VDD VSS sg13g2_FILL8
XSTDFILL78_608 VDD VSS sg13g2_FILL8
XSTDFILL78_616 VDD VSS sg13g2_FILL8
XSTDFILL78_624 VDD VSS sg13g2_FILL8
XSTDFILL78_632 VDD VSS sg13g2_FILL8
XSTDFILL78_640 VDD VSS sg13g2_FILL8
XSTDFILL78_648 VDD VSS sg13g2_FILL8
XSTDFILL78_656 VDD VSS sg13g2_FILL8
XSTDFILL78_664 VDD VSS sg13g2_FILL8
XSTDFILL78_672 VDD VSS sg13g2_FILL8
XSTDFILL78_680 VDD VSS sg13g2_FILL8
XSTDFILL78_688 VDD VSS sg13g2_FILL8
XSTDFILL78_696 VDD VSS sg13g2_FILL8
XSTDFILL78_704 VDD VSS sg13g2_FILL8
XSTDFILL78_712 VDD VSS sg13g2_FILL8
XSTDFILL78_720 VDD VSS sg13g2_FILL8
XSTDFILL78_728 VDD VSS sg13g2_FILL8
XSTDFILL78_736 VDD VSS sg13g2_FILL8
XSTDFILL78_744 VDD VSS sg13g2_FILL8
XSTDFILL78_752 VDD VSS sg13g2_FILL8
XSTDFILL78_760 VDD VSS sg13g2_FILL8
XSTDFILL78_768 VDD VSS sg13g2_FILL8
XSTDFILL78_776 VDD VSS sg13g2_FILL8
XSTDFILL78_784 VDD VSS sg13g2_FILL8
XSTDFILL78_792 VDD VSS sg13g2_FILL8
XSTDFILL78_800 VDD VSS sg13g2_FILL8
XSTDFILL78_808 VDD VSS sg13g2_FILL8
XSTDFILL78_816 VDD VSS sg13g2_FILL8
XSTDFILL78_824 VDD VSS sg13g2_FILL8
XSTDFILL78_832 VDD VSS sg13g2_FILL8
XSTDFILL78_840 VDD VSS sg13g2_FILL8
XSTDFILL78_848 VDD VSS sg13g2_FILL8
XSTDFILL78_856 VDD VSS sg13g2_FILL8
XSTDFILL78_864 VDD VSS sg13g2_FILL8
XSTDFILL78_872 VDD VSS sg13g2_FILL8
XSTDFILL78_880 VDD VSS sg13g2_FILL8
XSTDFILL78_888 VDD VSS sg13g2_FILL8
XSTDFILL78_896 VDD VSS sg13g2_FILL8
XSTDFILL78_904 VDD VSS sg13g2_FILL8
XSTDFILL78_912 VDD VSS sg13g2_FILL8
XSTDFILL78_920 VDD VSS sg13g2_FILL8
XSTDFILL78_928 VDD VSS sg13g2_FILL8
XSTDFILL78_936 VDD VSS sg13g2_FILL8
XSTDFILL78_944 VDD VSS sg13g2_FILL8
XSTDFILL78_952 VDD VSS sg13g2_FILL8
XSTDFILL78_960 VDD VSS sg13g2_FILL8
XSTDFILL78_968 VDD VSS sg13g2_FILL8
XSTDFILL78_976 VDD VSS sg13g2_FILL8
XSTDFILL78_984 VDD VSS sg13g2_FILL8
XSTDFILL78_992 VDD VSS sg13g2_FILL8
XSTDFILL78_1000 VDD VSS sg13g2_FILL8
XSTDFILL78_1008 VDD VSS sg13g2_FILL8
XSTDFILL78_1016 VDD VSS sg13g2_FILL8
XSTDFILL78_1024 VDD VSS sg13g2_FILL8
XSTDFILL78_1032 VDD VSS sg13g2_FILL8
XSTDFILL78_1040 VDD VSS sg13g2_FILL8
XSTDFILL78_1048 VDD VSS sg13g2_FILL8
XSTDFILL78_1056 VDD VSS sg13g2_FILL8
XSTDFILL78_1064 VDD VSS sg13g2_FILL8
XSTDFILL78_1072 VDD VSS sg13g2_FILL8
XSTDFILL78_1080 VDD VSS sg13g2_FILL8
XSTDFILL78_1088 VDD VSS sg13g2_FILL8
XSTDFILL78_1096 VDD VSS sg13g2_FILL8
XSTDFILL78_1104 VDD VSS sg13g2_FILL8
XSTDFILL78_1112 VDD VSS sg13g2_FILL8
XSTDFILL78_1120 VDD VSS sg13g2_FILL8
XSTDFILL78_1128 VDD VSS sg13g2_FILL8
XSTDFILL78_1136 VDD VSS sg13g2_FILL8
XSTDFILL78_1144 VDD VSS sg13g2_FILL8
XSTDFILL78_1152 VDD VSS sg13g2_FILL8
XSTDFILL78_1160 VDD VSS sg13g2_FILL8
XSTDFILL78_1168 VDD VSS sg13g2_FILL8
XSTDFILL78_1176 VDD VSS sg13g2_FILL8
XSTDFILL78_1184 VDD VSS sg13g2_FILL8
XSTDFILL78_1192 VDD VSS sg13g2_FILL8
XSTDFILL78_1200 VDD VSS sg13g2_FILL8
XSTDFILL78_1208 VDD VSS sg13g2_FILL8
XSTDFILL78_1216 VDD VSS sg13g2_FILL8
XSTDFILL78_1224 VDD VSS sg13g2_FILL8
XSTDFILL78_1232 VDD VSS sg13g2_FILL8
XSTDFILL78_1240 VDD VSS sg13g2_FILL8
XSTDFILL78_1248 VDD VSS sg13g2_FILL8
XSTDFILL78_1256 VDD VSS sg13g2_FILL8
XSTDFILL78_1264 VDD VSS sg13g2_FILL8
XSTDFILL78_1272 VDD VSS sg13g2_FILL8
XSTDFILL78_1280 VDD VSS sg13g2_FILL8
XSTDFILL78_1288 VDD VSS sg13g2_FILL8
XSTDFILL78_1296 VDD VSS sg13g2_FILL8
XSTDFILL78_1304 VDD VSS sg13g2_FILL8
XSTDFILL78_1312 VDD VSS sg13g2_FILL8
XSTDFILL78_1320 VDD VSS sg13g2_FILL8
XSTDFILL78_1328 VDD VSS sg13g2_FILL8
XSTDFILL78_1336 VDD VSS sg13g2_FILL8
XSTDFILL78_1344 VDD VSS sg13g2_FILL8
XSTDFILL78_1352 VDD VSS sg13g2_FILL8
XSTDFILL78_1360 VDD VSS sg13g2_FILL8
XSTDFILL78_1368 VDD VSS sg13g2_FILL8
XSTDFILL78_1376 VDD VSS sg13g2_FILL8
XSTDFILL78_1384 VDD VSS sg13g2_FILL8
XSTDFILL78_1392 VDD VSS sg13g2_FILL8
XSTDFILL78_1400 VDD VSS sg13g2_FILL8
XSTDFILL78_1408 VDD VSS sg13g2_FILL8
XSTDFILL78_1416 VDD VSS sg13g2_FILL8
XSTDFILL78_1424 VDD VSS sg13g2_FILL8
XSTDFILL78_1432 VDD VSS sg13g2_FILL8
XSTDFILL78_1440 VDD VSS sg13g2_FILL8
XSTDFILL78_1448 VDD VSS sg13g2_FILL8
XSTDFILL78_1456 VDD VSS sg13g2_FILL8
XSTDFILL78_1464 VDD VSS sg13g2_FILL8
XSTDFILL78_1472 VDD VSS sg13g2_FILL8
XSTDFILL78_1480 VDD VSS sg13g2_FILL8
XSTDFILL78_1488 VDD VSS sg13g2_FILL8
XSTDFILL78_1496 VDD VSS sg13g2_FILL8
XSTDFILL78_1504 VDD VSS sg13g2_FILL8
XSTDFILL78_1512 VDD VSS sg13g2_FILL8
XSTDFILL78_1520 VDD VSS sg13g2_FILL8
XSTDFILL78_1528 VDD VSS sg13g2_FILL2
XSTDFILL78_1530 VDD VSS sg13g2_FILL1
XSTDFILL79_0 VDD VSS sg13g2_FILL8
XSTDFILL79_8 VDD VSS sg13g2_FILL8
XSTDFILL79_16 VDD VSS sg13g2_FILL8
XSTDFILL79_24 VDD VSS sg13g2_FILL8
XSTDFILL79_32 VDD VSS sg13g2_FILL8
XSTDFILL79_40 VDD VSS sg13g2_FILL8
XSTDFILL79_48 VDD VSS sg13g2_FILL8
XSTDFILL79_56 VDD VSS sg13g2_FILL8
XSTDFILL79_64 VDD VSS sg13g2_FILL8
XSTDFILL79_72 VDD VSS sg13g2_FILL8
XSTDFILL79_80 VDD VSS sg13g2_FILL8
XSTDFILL79_88 VDD VSS sg13g2_FILL8
XSTDFILL79_96 VDD VSS sg13g2_FILL8
XSTDFILL79_104 VDD VSS sg13g2_FILL8
XSTDFILL79_112 VDD VSS sg13g2_FILL8
XSTDFILL79_120 VDD VSS sg13g2_FILL8
XSTDFILL79_128 VDD VSS sg13g2_FILL8
XSTDFILL79_136 VDD VSS sg13g2_FILL8
XSTDFILL79_144 VDD VSS sg13g2_FILL8
XSTDFILL79_152 VDD VSS sg13g2_FILL8
XSTDFILL79_160 VDD VSS sg13g2_FILL8
XSTDFILL79_168 VDD VSS sg13g2_FILL8
XSTDFILL79_176 VDD VSS sg13g2_FILL8
XSTDFILL79_184 VDD VSS sg13g2_FILL8
XSTDFILL79_192 VDD VSS sg13g2_FILL8
XSTDFILL79_200 VDD VSS sg13g2_FILL8
XSTDFILL79_208 VDD VSS sg13g2_FILL8
XSTDFILL79_216 VDD VSS sg13g2_FILL8
XSTDFILL79_224 VDD VSS sg13g2_FILL8
XSTDFILL79_232 VDD VSS sg13g2_FILL8
XSTDFILL79_240 VDD VSS sg13g2_FILL8
XSTDFILL79_248 VDD VSS sg13g2_FILL8
XSTDFILL79_256 VDD VSS sg13g2_FILL8
XSTDFILL79_264 VDD VSS sg13g2_FILL8
XSTDFILL79_272 VDD VSS sg13g2_FILL8
XSTDFILL79_280 VDD VSS sg13g2_FILL8
XSTDFILL79_288 VDD VSS sg13g2_FILL8
XSTDFILL79_296 VDD VSS sg13g2_FILL8
XSTDFILL79_304 VDD VSS sg13g2_FILL8
XSTDFILL79_312 VDD VSS sg13g2_FILL8
XSTDFILL79_320 VDD VSS sg13g2_FILL8
XSTDFILL79_328 VDD VSS sg13g2_FILL8
XSTDFILL79_336 VDD VSS sg13g2_FILL8
XSTDFILL79_344 VDD VSS sg13g2_FILL8
XSTDFILL79_352 VDD VSS sg13g2_FILL8
XSTDFILL79_360 VDD VSS sg13g2_FILL8
XSTDFILL79_368 VDD VSS sg13g2_FILL8
XSTDFILL79_376 VDD VSS sg13g2_FILL8
XSTDFILL79_384 VDD VSS sg13g2_FILL8
XSTDFILL79_392 VDD VSS sg13g2_FILL8
XSTDFILL79_400 VDD VSS sg13g2_FILL8
XSTDFILL79_408 VDD VSS sg13g2_FILL8
XSTDFILL79_416 VDD VSS sg13g2_FILL8
XSTDFILL79_424 VDD VSS sg13g2_FILL8
XSTDFILL79_432 VDD VSS sg13g2_FILL8
XSTDFILL79_440 VDD VSS sg13g2_FILL8
XSTDFILL79_448 VDD VSS sg13g2_FILL8
XSTDFILL79_456 VDD VSS sg13g2_FILL8
XSTDFILL79_464 VDD VSS sg13g2_FILL8
XSTDFILL79_472 VDD VSS sg13g2_FILL8
XSTDFILL79_480 VDD VSS sg13g2_FILL8
XSTDFILL79_488 VDD VSS sg13g2_FILL8
XSTDFILL79_496 VDD VSS sg13g2_FILL8
XSTDFILL79_504 VDD VSS sg13g2_FILL8
XSTDFILL79_512 VDD VSS sg13g2_FILL8
XSTDFILL79_520 VDD VSS sg13g2_FILL8
XSTDFILL79_528 VDD VSS sg13g2_FILL8
XSTDFILL79_536 VDD VSS sg13g2_FILL8
XSTDFILL79_544 VDD VSS sg13g2_FILL8
XSTDFILL79_552 VDD VSS sg13g2_FILL8
XSTDFILL79_560 VDD VSS sg13g2_FILL8
XSTDFILL79_568 VDD VSS sg13g2_FILL8
XSTDFILL79_576 VDD VSS sg13g2_FILL8
XSTDFILL79_584 VDD VSS sg13g2_FILL8
XSTDFILL79_592 VDD VSS sg13g2_FILL8
XSTDFILL79_600 VDD VSS sg13g2_FILL8
XSTDFILL79_608 VDD VSS sg13g2_FILL8
XSTDFILL79_616 VDD VSS sg13g2_FILL8
XSTDFILL79_624 VDD VSS sg13g2_FILL8
XSTDFILL79_632 VDD VSS sg13g2_FILL8
XSTDFILL79_640 VDD VSS sg13g2_FILL8
XSTDFILL79_648 VDD VSS sg13g2_FILL8
XSTDFILL79_656 VDD VSS sg13g2_FILL8
XSTDFILL79_664 VDD VSS sg13g2_FILL8
XSTDFILL79_672 VDD VSS sg13g2_FILL8
XSTDFILL79_680 VDD VSS sg13g2_FILL8
XSTDFILL79_688 VDD VSS sg13g2_FILL8
XSTDFILL79_696 VDD VSS sg13g2_FILL8
XSTDFILL79_704 VDD VSS sg13g2_FILL8
XSTDFILL79_712 VDD VSS sg13g2_FILL8
XSTDFILL79_720 VDD VSS sg13g2_FILL8
XSTDFILL79_728 VDD VSS sg13g2_FILL8
XSTDFILL79_736 VDD VSS sg13g2_FILL8
XSTDFILL79_744 VDD VSS sg13g2_FILL8
XSTDFILL79_752 VDD VSS sg13g2_FILL8
XSTDFILL79_760 VDD VSS sg13g2_FILL8
XSTDFILL79_768 VDD VSS sg13g2_FILL8
XSTDFILL79_776 VDD VSS sg13g2_FILL8
XSTDFILL79_784 VDD VSS sg13g2_FILL8
XSTDFILL79_792 VDD VSS sg13g2_FILL8
XSTDFILL79_800 VDD VSS sg13g2_FILL8
XSTDFILL79_808 VDD VSS sg13g2_FILL8
XSTDFILL79_816 VDD VSS sg13g2_FILL8
XSTDFILL79_824 VDD VSS sg13g2_FILL8
XSTDFILL79_832 VDD VSS sg13g2_FILL8
XSTDFILL79_840 VDD VSS sg13g2_FILL8
XSTDFILL79_848 VDD VSS sg13g2_FILL8
XSTDFILL79_856 VDD VSS sg13g2_FILL8
XSTDFILL79_864 VDD VSS sg13g2_FILL8
XSTDFILL79_872 VDD VSS sg13g2_FILL8
XSTDFILL79_880 VDD VSS sg13g2_FILL8
XSTDFILL79_888 VDD VSS sg13g2_FILL8
XSTDFILL79_896 VDD VSS sg13g2_FILL8
XSTDFILL79_904 VDD VSS sg13g2_FILL8
XSTDFILL79_912 VDD VSS sg13g2_FILL8
XSTDFILL79_920 VDD VSS sg13g2_FILL8
XSTDFILL79_928 VDD VSS sg13g2_FILL8
XSTDFILL79_936 VDD VSS sg13g2_FILL8
XSTDFILL79_944 VDD VSS sg13g2_FILL8
XSTDFILL79_952 VDD VSS sg13g2_FILL8
XSTDFILL79_960 VDD VSS sg13g2_FILL8
XSTDFILL79_968 VDD VSS sg13g2_FILL8
XSTDFILL79_976 VDD VSS sg13g2_FILL8
XSTDFILL79_984 VDD VSS sg13g2_FILL8
XSTDFILL79_992 VDD VSS sg13g2_FILL8
XSTDFILL79_1000 VDD VSS sg13g2_FILL8
XSTDFILL79_1008 VDD VSS sg13g2_FILL8
XSTDFILL79_1016 VDD VSS sg13g2_FILL8
XSTDFILL79_1024 VDD VSS sg13g2_FILL8
XSTDFILL79_1032 VDD VSS sg13g2_FILL8
XSTDFILL79_1040 VDD VSS sg13g2_FILL8
XSTDFILL79_1048 VDD VSS sg13g2_FILL8
XSTDFILL79_1056 VDD VSS sg13g2_FILL8
XSTDFILL79_1064 VDD VSS sg13g2_FILL8
XSTDFILL79_1072 VDD VSS sg13g2_FILL8
XSTDFILL79_1080 VDD VSS sg13g2_FILL8
XSTDFILL79_1088 VDD VSS sg13g2_FILL8
XSTDFILL79_1096 VDD VSS sg13g2_FILL8
XSTDFILL79_1104 VDD VSS sg13g2_FILL8
XSTDFILL79_1112 VDD VSS sg13g2_FILL8
XSTDFILL79_1120 VDD VSS sg13g2_FILL8
XSTDFILL79_1128 VDD VSS sg13g2_FILL8
XSTDFILL79_1136 VDD VSS sg13g2_FILL8
XSTDFILL79_1144 VDD VSS sg13g2_FILL8
XSTDFILL79_1152 VDD VSS sg13g2_FILL8
XSTDFILL79_1160 VDD VSS sg13g2_FILL8
XSTDFILL79_1168 VDD VSS sg13g2_FILL8
XSTDFILL79_1176 VDD VSS sg13g2_FILL8
XSTDFILL79_1184 VDD VSS sg13g2_FILL8
XSTDFILL79_1192 VDD VSS sg13g2_FILL8
XSTDFILL79_1200 VDD VSS sg13g2_FILL8
XSTDFILL79_1208 VDD VSS sg13g2_FILL8
XSTDFILL79_1216 VDD VSS sg13g2_FILL8
XSTDFILL79_1224 VDD VSS sg13g2_FILL8
XSTDFILL79_1232 VDD VSS sg13g2_FILL8
XSTDFILL79_1240 VDD VSS sg13g2_FILL8
XSTDFILL79_1248 VDD VSS sg13g2_FILL8
XSTDFILL79_1256 VDD VSS sg13g2_FILL8
XSTDFILL79_1264 VDD VSS sg13g2_FILL8
XSTDFILL79_1272 VDD VSS sg13g2_FILL8
XSTDFILL79_1280 VDD VSS sg13g2_FILL8
XSTDFILL79_1288 VDD VSS sg13g2_FILL8
XSTDFILL79_1296 VDD VSS sg13g2_FILL8
XSTDFILL79_1304 VDD VSS sg13g2_FILL8
XSTDFILL79_1312 VDD VSS sg13g2_FILL8
XSTDFILL79_1320 VDD VSS sg13g2_FILL8
XSTDFILL79_1328 VDD VSS sg13g2_FILL8
XSTDFILL79_1336 VDD VSS sg13g2_FILL8
XSTDFILL79_1344 VDD VSS sg13g2_FILL8
XSTDFILL79_1352 VDD VSS sg13g2_FILL8
XSTDFILL79_1360 VDD VSS sg13g2_FILL8
XSTDFILL79_1368 VDD VSS sg13g2_FILL8
XSTDFILL79_1376 VDD VSS sg13g2_FILL8
XSTDFILL79_1384 VDD VSS sg13g2_FILL8
XSTDFILL79_1392 VDD VSS sg13g2_FILL8
XSTDFILL79_1400 VDD VSS sg13g2_FILL8
XSTDFILL79_1408 VDD VSS sg13g2_FILL8
XSTDFILL79_1416 VDD VSS sg13g2_FILL8
XSTDFILL79_1424 VDD VSS sg13g2_FILL8
XSTDFILL79_1432 VDD VSS sg13g2_FILL8
XSTDFILL79_1440 VDD VSS sg13g2_FILL8
XSTDFILL79_1448 VDD VSS sg13g2_FILL8
XSTDFILL79_1456 VDD VSS sg13g2_FILL8
XSTDFILL79_1464 VDD VSS sg13g2_FILL8
XSTDFILL79_1472 VDD VSS sg13g2_FILL8
XSTDFILL79_1480 VDD VSS sg13g2_FILL8
XSTDFILL79_1488 VDD VSS sg13g2_FILL8
XSTDFILL79_1496 VDD VSS sg13g2_FILL8
XSTDFILL79_1504 VDD VSS sg13g2_FILL8
XSTDFILL79_1512 VDD VSS sg13g2_FILL8
XSTDFILL79_1520 VDD VSS sg13g2_FILL8
XSTDFILL79_1528 VDD VSS sg13g2_FILL2
XSTDFILL79_1530 VDD VSS sg13g2_FILL1
XSTDFILL80_0 VDD VSS sg13g2_FILL8
XSTDFILL80_8 VDD VSS sg13g2_FILL8
XSTDFILL80_16 VDD VSS sg13g2_FILL8
XSTDFILL80_24 VDD VSS sg13g2_FILL8
XSTDFILL80_32 VDD VSS sg13g2_FILL8
XSTDFILL80_40 VDD VSS sg13g2_FILL8
XSTDFILL80_48 VDD VSS sg13g2_FILL8
XSTDFILL80_56 VDD VSS sg13g2_FILL8
XSTDFILL80_64 VDD VSS sg13g2_FILL8
XSTDFILL80_72 VDD VSS sg13g2_FILL8
XSTDFILL80_80 VDD VSS sg13g2_FILL8
XSTDFILL80_88 VDD VSS sg13g2_FILL8
XSTDFILL80_96 VDD VSS sg13g2_FILL8
XSTDFILL80_104 VDD VSS sg13g2_FILL8
XSTDFILL80_112 VDD VSS sg13g2_FILL8
XSTDFILL80_120 VDD VSS sg13g2_FILL8
XSTDFILL80_128 VDD VSS sg13g2_FILL8
XSTDFILL80_136 VDD VSS sg13g2_FILL8
XSTDFILL80_144 VDD VSS sg13g2_FILL8
XSTDFILL80_152 VDD VSS sg13g2_FILL8
XSTDFILL80_160 VDD VSS sg13g2_FILL8
XSTDFILL80_168 VDD VSS sg13g2_FILL8
XSTDFILL80_176 VDD VSS sg13g2_FILL8
XSTDFILL80_184 VDD VSS sg13g2_FILL8
XSTDFILL80_192 VDD VSS sg13g2_FILL8
XSTDFILL80_200 VDD VSS sg13g2_FILL8
XSTDFILL80_208 VDD VSS sg13g2_FILL8
XSTDFILL80_216 VDD VSS sg13g2_FILL8
XSTDFILL80_224 VDD VSS sg13g2_FILL8
XSTDFILL80_232 VDD VSS sg13g2_FILL8
XSTDFILL80_240 VDD VSS sg13g2_FILL8
XSTDFILL80_248 VDD VSS sg13g2_FILL8
XSTDFILL80_256 VDD VSS sg13g2_FILL8
XSTDFILL80_264 VDD VSS sg13g2_FILL8
XSTDFILL80_272 VDD VSS sg13g2_FILL8
XSTDFILL80_280 VDD VSS sg13g2_FILL8
XSTDFILL80_288 VDD VSS sg13g2_FILL8
XSTDFILL80_296 VDD VSS sg13g2_FILL8
XSTDFILL80_304 VDD VSS sg13g2_FILL8
XSTDFILL80_312 VDD VSS sg13g2_FILL8
XSTDFILL80_320 VDD VSS sg13g2_FILL8
XSTDFILL80_328 VDD VSS sg13g2_FILL8
XSTDFILL80_336 VDD VSS sg13g2_FILL8
XSTDFILL80_344 VDD VSS sg13g2_FILL8
XSTDFILL80_352 VDD VSS sg13g2_FILL8
XSTDFILL80_360 VDD VSS sg13g2_FILL8
XSTDFILL80_368 VDD VSS sg13g2_FILL8
XSTDFILL80_376 VDD VSS sg13g2_FILL8
XSTDFILL80_384 VDD VSS sg13g2_FILL8
XSTDFILL80_392 VDD VSS sg13g2_FILL8
XSTDFILL80_400 VDD VSS sg13g2_FILL8
XSTDFILL80_408 VDD VSS sg13g2_FILL8
XSTDFILL80_416 VDD VSS sg13g2_FILL8
XSTDFILL80_424 VDD VSS sg13g2_FILL8
XSTDFILL80_432 VDD VSS sg13g2_FILL8
XSTDFILL80_440 VDD VSS sg13g2_FILL8
XSTDFILL80_448 VDD VSS sg13g2_FILL8
XSTDFILL80_456 VDD VSS sg13g2_FILL8
XSTDFILL80_464 VDD VSS sg13g2_FILL8
XSTDFILL80_472 VDD VSS sg13g2_FILL8
XSTDFILL80_480 VDD VSS sg13g2_FILL8
XSTDFILL80_488 VDD VSS sg13g2_FILL8
XSTDFILL80_496 VDD VSS sg13g2_FILL8
XSTDFILL80_504 VDD VSS sg13g2_FILL8
XSTDFILL80_512 VDD VSS sg13g2_FILL8
XSTDFILL80_520 VDD VSS sg13g2_FILL8
XSTDFILL80_528 VDD VSS sg13g2_FILL8
XSTDFILL80_536 VDD VSS sg13g2_FILL8
XSTDFILL80_544 VDD VSS sg13g2_FILL8
XSTDFILL80_552 VDD VSS sg13g2_FILL8
XSTDFILL80_560 VDD VSS sg13g2_FILL8
XSTDFILL80_568 VDD VSS sg13g2_FILL8
XSTDFILL80_576 VDD VSS sg13g2_FILL8
XSTDFILL80_584 VDD VSS sg13g2_FILL8
XSTDFILL80_592 VDD VSS sg13g2_FILL8
XSTDFILL80_600 VDD VSS sg13g2_FILL8
XSTDFILL80_608 VDD VSS sg13g2_FILL8
XSTDFILL80_616 VDD VSS sg13g2_FILL8
XSTDFILL80_624 VDD VSS sg13g2_FILL8
XSTDFILL80_632 VDD VSS sg13g2_FILL8
XSTDFILL80_640 VDD VSS sg13g2_FILL8
XSTDFILL80_648 VDD VSS sg13g2_FILL8
XSTDFILL80_656 VDD VSS sg13g2_FILL8
XSTDFILL80_664 VDD VSS sg13g2_FILL8
XSTDFILL80_672 VDD VSS sg13g2_FILL8
XSTDFILL80_680 VDD VSS sg13g2_FILL8
XSTDFILL80_688 VDD VSS sg13g2_FILL8
XSTDFILL80_696 VDD VSS sg13g2_FILL8
XSTDFILL80_704 VDD VSS sg13g2_FILL8
XSTDFILL80_712 VDD VSS sg13g2_FILL8
XSTDFILL80_720 VDD VSS sg13g2_FILL8
XSTDFILL80_728 VDD VSS sg13g2_FILL8
XSTDFILL80_736 VDD VSS sg13g2_FILL8
XSTDFILL80_744 VDD VSS sg13g2_FILL8
XSTDFILL80_752 VDD VSS sg13g2_FILL8
XSTDFILL80_760 VDD VSS sg13g2_FILL8
XSTDFILL80_768 VDD VSS sg13g2_FILL8
XSTDFILL80_776 VDD VSS sg13g2_FILL8
XSTDFILL80_784 VDD VSS sg13g2_FILL8
XSTDFILL80_792 VDD VSS sg13g2_FILL8
XSTDFILL80_800 VDD VSS sg13g2_FILL8
XSTDFILL80_808 VDD VSS sg13g2_FILL8
XSTDFILL80_816 VDD VSS sg13g2_FILL8
XSTDFILL80_824 VDD VSS sg13g2_FILL8
XSTDFILL80_832 VDD VSS sg13g2_FILL8
XSTDFILL80_840 VDD VSS sg13g2_FILL8
XSTDFILL80_848 VDD VSS sg13g2_FILL8
XSTDFILL80_856 VDD VSS sg13g2_FILL8
XSTDFILL80_864 VDD VSS sg13g2_FILL8
XSTDFILL80_872 VDD VSS sg13g2_FILL8
XSTDFILL80_880 VDD VSS sg13g2_FILL8
XSTDFILL80_888 VDD VSS sg13g2_FILL8
XSTDFILL80_896 VDD VSS sg13g2_FILL8
XSTDFILL80_904 VDD VSS sg13g2_FILL8
XSTDFILL80_912 VDD VSS sg13g2_FILL8
XSTDFILL80_920 VDD VSS sg13g2_FILL8
XSTDFILL80_928 VDD VSS sg13g2_FILL8
XSTDFILL80_936 VDD VSS sg13g2_FILL8
XSTDFILL80_944 VDD VSS sg13g2_FILL8
XSTDFILL80_952 VDD VSS sg13g2_FILL8
XSTDFILL80_960 VDD VSS sg13g2_FILL8
XSTDFILL80_968 VDD VSS sg13g2_FILL8
XSTDFILL80_976 VDD VSS sg13g2_FILL8
XSTDFILL80_984 VDD VSS sg13g2_FILL8
XSTDFILL80_992 VDD VSS sg13g2_FILL8
XSTDFILL80_1000 VDD VSS sg13g2_FILL8
XSTDFILL80_1008 VDD VSS sg13g2_FILL8
XSTDFILL80_1016 VDD VSS sg13g2_FILL8
XSTDFILL80_1024 VDD VSS sg13g2_FILL8
XSTDFILL80_1032 VDD VSS sg13g2_FILL8
XSTDFILL80_1040 VDD VSS sg13g2_FILL8
XSTDFILL80_1048 VDD VSS sg13g2_FILL8
XSTDFILL80_1056 VDD VSS sg13g2_FILL8
XSTDFILL80_1064 VDD VSS sg13g2_FILL8
XSTDFILL80_1072 VDD VSS sg13g2_FILL8
XSTDFILL80_1080 VDD VSS sg13g2_FILL8
XSTDFILL80_1088 VDD VSS sg13g2_FILL8
XSTDFILL80_1096 VDD VSS sg13g2_FILL8
XSTDFILL80_1104 VDD VSS sg13g2_FILL8
XSTDFILL80_1112 VDD VSS sg13g2_FILL8
XSTDFILL80_1120 VDD VSS sg13g2_FILL8
XSTDFILL80_1128 VDD VSS sg13g2_FILL8
XSTDFILL80_1136 VDD VSS sg13g2_FILL8
XSTDFILL80_1144 VDD VSS sg13g2_FILL8
XSTDFILL80_1152 VDD VSS sg13g2_FILL8
XSTDFILL80_1160 VDD VSS sg13g2_FILL8
XSTDFILL80_1168 VDD VSS sg13g2_FILL8
XSTDFILL80_1176 VDD VSS sg13g2_FILL8
XSTDFILL80_1184 VDD VSS sg13g2_FILL8
XSTDFILL80_1192 VDD VSS sg13g2_FILL8
XSTDFILL80_1200 VDD VSS sg13g2_FILL8
XSTDFILL80_1208 VDD VSS sg13g2_FILL8
XSTDFILL80_1216 VDD VSS sg13g2_FILL8
XSTDFILL80_1224 VDD VSS sg13g2_FILL8
XSTDFILL80_1232 VDD VSS sg13g2_FILL8
XSTDFILL80_1240 VDD VSS sg13g2_FILL8
XSTDFILL80_1248 VDD VSS sg13g2_FILL8
XSTDFILL80_1256 VDD VSS sg13g2_FILL8
XSTDFILL80_1264 VDD VSS sg13g2_FILL8
XSTDFILL80_1272 VDD VSS sg13g2_FILL8
XSTDFILL80_1280 VDD VSS sg13g2_FILL8
XSTDFILL80_1288 VDD VSS sg13g2_FILL8
XSTDFILL80_1296 VDD VSS sg13g2_FILL8
XSTDFILL80_1304 VDD VSS sg13g2_FILL8
XSTDFILL80_1312 VDD VSS sg13g2_FILL8
XSTDFILL80_1320 VDD VSS sg13g2_FILL8
XSTDFILL80_1328 VDD VSS sg13g2_FILL8
XSTDFILL80_1336 VDD VSS sg13g2_FILL8
XSTDFILL80_1344 VDD VSS sg13g2_FILL8
XSTDFILL80_1352 VDD VSS sg13g2_FILL8
XSTDFILL80_1360 VDD VSS sg13g2_FILL8
XSTDFILL80_1368 VDD VSS sg13g2_FILL8
XSTDFILL80_1376 VDD VSS sg13g2_FILL8
XSTDFILL80_1384 VDD VSS sg13g2_FILL8
XSTDFILL80_1392 VDD VSS sg13g2_FILL8
XSTDFILL80_1400 VDD VSS sg13g2_FILL8
XSTDFILL80_1408 VDD VSS sg13g2_FILL8
XSTDFILL80_1416 VDD VSS sg13g2_FILL8
XSTDFILL80_1424 VDD VSS sg13g2_FILL8
XSTDFILL80_1432 VDD VSS sg13g2_FILL8
XSTDFILL80_1440 VDD VSS sg13g2_FILL8
XSTDFILL80_1448 VDD VSS sg13g2_FILL8
XSTDFILL80_1456 VDD VSS sg13g2_FILL8
XSTDFILL80_1464 VDD VSS sg13g2_FILL8
XSTDFILL80_1472 VDD VSS sg13g2_FILL8
XSTDFILL80_1480 VDD VSS sg13g2_FILL8
XSTDFILL80_1488 VDD VSS sg13g2_FILL8
XSTDFILL80_1496 VDD VSS sg13g2_FILL8
XSTDFILL80_1504 VDD VSS sg13g2_FILL8
XSTDFILL80_1512 VDD VSS sg13g2_FILL8
XSTDFILL80_1520 VDD VSS sg13g2_FILL8
XSTDFILL80_1528 VDD VSS sg13g2_FILL2
XSTDFILL80_1530 VDD VSS sg13g2_FILL1
XSTDFILL81_0 VDD VSS sg13g2_FILL8
XSTDFILL81_8 VDD VSS sg13g2_FILL8
XSTDFILL81_16 VDD VSS sg13g2_FILL8
XSTDFILL81_24 VDD VSS sg13g2_FILL8
XSTDFILL81_32 VDD VSS sg13g2_FILL8
XSTDFILL81_40 VDD VSS sg13g2_FILL8
XSTDFILL81_48 VDD VSS sg13g2_FILL8
XSTDFILL81_56 VDD VSS sg13g2_FILL8
XSTDFILL81_64 VDD VSS sg13g2_FILL8
XSTDFILL81_72 VDD VSS sg13g2_FILL8
XSTDFILL81_80 VDD VSS sg13g2_FILL8
XSTDFILL81_88 VDD VSS sg13g2_FILL8
XSTDFILL81_96 VDD VSS sg13g2_FILL8
XSTDFILL81_104 VDD VSS sg13g2_FILL8
XSTDFILL81_112 VDD VSS sg13g2_FILL8
XSTDFILL81_120 VDD VSS sg13g2_FILL8
XSTDFILL81_128 VDD VSS sg13g2_FILL8
XSTDFILL81_136 VDD VSS sg13g2_FILL8
XSTDFILL81_144 VDD VSS sg13g2_FILL8
XSTDFILL81_152 VDD VSS sg13g2_FILL8
XSTDFILL81_160 VDD VSS sg13g2_FILL8
XSTDFILL81_168 VDD VSS sg13g2_FILL8
XSTDFILL81_176 VDD VSS sg13g2_FILL8
XSTDFILL81_184 VDD VSS sg13g2_FILL8
XSTDFILL81_192 VDD VSS sg13g2_FILL8
XSTDFILL81_200 VDD VSS sg13g2_FILL8
XSTDFILL81_208 VDD VSS sg13g2_FILL8
XSTDFILL81_216 VDD VSS sg13g2_FILL8
XSTDFILL81_224 VDD VSS sg13g2_FILL8
XSTDFILL81_232 VDD VSS sg13g2_FILL8
XSTDFILL81_240 VDD VSS sg13g2_FILL8
XSTDFILL81_248 VDD VSS sg13g2_FILL8
XSTDFILL81_256 VDD VSS sg13g2_FILL8
XSTDFILL81_264 VDD VSS sg13g2_FILL8
XSTDFILL81_272 VDD VSS sg13g2_FILL8
XSTDFILL81_280 VDD VSS sg13g2_FILL8
XSTDFILL81_288 VDD VSS sg13g2_FILL8
XSTDFILL81_296 VDD VSS sg13g2_FILL8
XSTDFILL81_304 VDD VSS sg13g2_FILL8
XSTDFILL81_312 VDD VSS sg13g2_FILL8
XSTDFILL81_320 VDD VSS sg13g2_FILL8
XSTDFILL81_328 VDD VSS sg13g2_FILL8
XSTDFILL81_336 VDD VSS sg13g2_FILL8
XSTDFILL81_344 VDD VSS sg13g2_FILL8
XSTDFILL81_352 VDD VSS sg13g2_FILL8
XSTDFILL81_360 VDD VSS sg13g2_FILL8
XSTDFILL81_368 VDD VSS sg13g2_FILL8
XSTDFILL81_376 VDD VSS sg13g2_FILL8
XSTDFILL81_384 VDD VSS sg13g2_FILL8
XSTDFILL81_392 VDD VSS sg13g2_FILL8
XSTDFILL81_400 VDD VSS sg13g2_FILL8
XSTDFILL81_408 VDD VSS sg13g2_FILL8
XSTDFILL81_416 VDD VSS sg13g2_FILL8
XSTDFILL81_424 VDD VSS sg13g2_FILL8
XSTDFILL81_432 VDD VSS sg13g2_FILL8
XSTDFILL81_440 VDD VSS sg13g2_FILL8
XSTDFILL81_448 VDD VSS sg13g2_FILL8
XSTDFILL81_456 VDD VSS sg13g2_FILL8
XSTDFILL81_464 VDD VSS sg13g2_FILL8
XSTDFILL81_472 VDD VSS sg13g2_FILL8
XSTDFILL81_480 VDD VSS sg13g2_FILL8
XSTDFILL81_488 VDD VSS sg13g2_FILL8
XSTDFILL81_496 VDD VSS sg13g2_FILL8
XSTDFILL81_504 VDD VSS sg13g2_FILL8
XSTDFILL81_512 VDD VSS sg13g2_FILL8
XSTDFILL81_520 VDD VSS sg13g2_FILL8
XSTDFILL81_528 VDD VSS sg13g2_FILL8
XSTDFILL81_536 VDD VSS sg13g2_FILL8
XSTDFILL81_544 VDD VSS sg13g2_FILL8
XSTDFILL81_552 VDD VSS sg13g2_FILL8
XSTDFILL81_560 VDD VSS sg13g2_FILL8
XSTDFILL81_568 VDD VSS sg13g2_FILL8
XSTDFILL81_576 VDD VSS sg13g2_FILL8
XSTDFILL81_584 VDD VSS sg13g2_FILL8
XSTDFILL81_592 VDD VSS sg13g2_FILL8
XSTDFILL81_600 VDD VSS sg13g2_FILL8
XSTDFILL81_608 VDD VSS sg13g2_FILL8
XSTDFILL81_616 VDD VSS sg13g2_FILL8
XSTDFILL81_624 VDD VSS sg13g2_FILL8
XSTDFILL81_632 VDD VSS sg13g2_FILL8
XSTDFILL81_640 VDD VSS sg13g2_FILL8
XSTDFILL81_648 VDD VSS sg13g2_FILL8
XSTDFILL81_656 VDD VSS sg13g2_FILL8
XSTDFILL81_664 VDD VSS sg13g2_FILL8
XSTDFILL81_672 VDD VSS sg13g2_FILL8
XSTDFILL81_680 VDD VSS sg13g2_FILL8
XSTDFILL81_688 VDD VSS sg13g2_FILL8
XSTDFILL81_696 VDD VSS sg13g2_FILL8
XSTDFILL81_704 VDD VSS sg13g2_FILL8
XSTDFILL81_712 VDD VSS sg13g2_FILL8
XSTDFILL81_720 VDD VSS sg13g2_FILL8
XSTDFILL81_728 VDD VSS sg13g2_FILL8
XSTDFILL81_736 VDD VSS sg13g2_FILL8
XSTDFILL81_744 VDD VSS sg13g2_FILL8
XSTDFILL81_752 VDD VSS sg13g2_FILL8
XSTDFILL81_760 VDD VSS sg13g2_FILL8
XSTDFILL81_768 VDD VSS sg13g2_FILL8
XSTDFILL81_776 VDD VSS sg13g2_FILL8
XSTDFILL81_784 VDD VSS sg13g2_FILL8
XSTDFILL81_792 VDD VSS sg13g2_FILL8
XSTDFILL81_800 VDD VSS sg13g2_FILL8
XSTDFILL81_808 VDD VSS sg13g2_FILL8
XSTDFILL81_816 VDD VSS sg13g2_FILL8
XSTDFILL81_824 VDD VSS sg13g2_FILL8
XSTDFILL81_832 VDD VSS sg13g2_FILL8
XSTDFILL81_840 VDD VSS sg13g2_FILL8
XSTDFILL81_848 VDD VSS sg13g2_FILL8
XSTDFILL81_856 VDD VSS sg13g2_FILL8
XSTDFILL81_864 VDD VSS sg13g2_FILL8
XSTDFILL81_872 VDD VSS sg13g2_FILL8
XSTDFILL81_880 VDD VSS sg13g2_FILL8
XSTDFILL81_888 VDD VSS sg13g2_FILL8
XSTDFILL81_896 VDD VSS sg13g2_FILL8
XSTDFILL81_904 VDD VSS sg13g2_FILL8
XSTDFILL81_912 VDD VSS sg13g2_FILL8
XSTDFILL81_920 VDD VSS sg13g2_FILL8
XSTDFILL81_928 VDD VSS sg13g2_FILL8
XSTDFILL81_936 VDD VSS sg13g2_FILL8
XSTDFILL81_944 VDD VSS sg13g2_FILL8
XSTDFILL81_952 VDD VSS sg13g2_FILL8
XSTDFILL81_960 VDD VSS sg13g2_FILL8
XSTDFILL81_968 VDD VSS sg13g2_FILL8
XSTDFILL81_976 VDD VSS sg13g2_FILL8
XSTDFILL81_984 VDD VSS sg13g2_FILL8
XSTDFILL81_992 VDD VSS sg13g2_FILL8
XSTDFILL81_1000 VDD VSS sg13g2_FILL8
XSTDFILL81_1008 VDD VSS sg13g2_FILL8
XSTDFILL81_1016 VDD VSS sg13g2_FILL8
XSTDFILL81_1024 VDD VSS sg13g2_FILL8
XSTDFILL81_1032 VDD VSS sg13g2_FILL8
XSTDFILL81_1040 VDD VSS sg13g2_FILL8
XSTDFILL81_1048 VDD VSS sg13g2_FILL8
XSTDFILL81_1056 VDD VSS sg13g2_FILL8
XSTDFILL81_1064 VDD VSS sg13g2_FILL8
XSTDFILL81_1072 VDD VSS sg13g2_FILL8
XSTDFILL81_1080 VDD VSS sg13g2_FILL8
XSTDFILL81_1088 VDD VSS sg13g2_FILL8
XSTDFILL81_1096 VDD VSS sg13g2_FILL8
XSTDFILL81_1104 VDD VSS sg13g2_FILL8
XSTDFILL81_1112 VDD VSS sg13g2_FILL8
XSTDFILL81_1120 VDD VSS sg13g2_FILL8
XSTDFILL81_1128 VDD VSS sg13g2_FILL8
XSTDFILL81_1136 VDD VSS sg13g2_FILL8
XSTDFILL81_1144 VDD VSS sg13g2_FILL8
XSTDFILL81_1152 VDD VSS sg13g2_FILL8
XSTDFILL81_1160 VDD VSS sg13g2_FILL8
XSTDFILL81_1168 VDD VSS sg13g2_FILL8
XSTDFILL81_1176 VDD VSS sg13g2_FILL8
XSTDFILL81_1184 VDD VSS sg13g2_FILL8
XSTDFILL81_1192 VDD VSS sg13g2_FILL8
XSTDFILL81_1200 VDD VSS sg13g2_FILL8
XSTDFILL81_1208 VDD VSS sg13g2_FILL8
XSTDFILL81_1216 VDD VSS sg13g2_FILL8
XSTDFILL81_1224 VDD VSS sg13g2_FILL8
XSTDFILL81_1232 VDD VSS sg13g2_FILL8
XSTDFILL81_1240 VDD VSS sg13g2_FILL8
XSTDFILL81_1248 VDD VSS sg13g2_FILL8
XSTDFILL81_1256 VDD VSS sg13g2_FILL8
XSTDFILL81_1264 VDD VSS sg13g2_FILL8
XSTDFILL81_1272 VDD VSS sg13g2_FILL8
XSTDFILL81_1280 VDD VSS sg13g2_FILL8
XSTDFILL81_1288 VDD VSS sg13g2_FILL8
XSTDFILL81_1296 VDD VSS sg13g2_FILL8
XSTDFILL81_1304 VDD VSS sg13g2_FILL8
XSTDFILL81_1312 VDD VSS sg13g2_FILL8
XSTDFILL81_1320 VDD VSS sg13g2_FILL8
XSTDFILL81_1328 VDD VSS sg13g2_FILL8
XSTDFILL81_1336 VDD VSS sg13g2_FILL8
XSTDFILL81_1344 VDD VSS sg13g2_FILL8
XSTDFILL81_1352 VDD VSS sg13g2_FILL8
XSTDFILL81_1360 VDD VSS sg13g2_FILL8
XSTDFILL81_1368 VDD VSS sg13g2_FILL8
XSTDFILL81_1376 VDD VSS sg13g2_FILL8
XSTDFILL81_1384 VDD VSS sg13g2_FILL8
XSTDFILL81_1392 VDD VSS sg13g2_FILL8
XSTDFILL81_1400 VDD VSS sg13g2_FILL8
XSTDFILL81_1408 VDD VSS sg13g2_FILL8
XSTDFILL81_1416 VDD VSS sg13g2_FILL8
XSTDFILL81_1424 VDD VSS sg13g2_FILL8
XSTDFILL81_1432 VDD VSS sg13g2_FILL8
XSTDFILL81_1440 VDD VSS sg13g2_FILL8
XSTDFILL81_1448 VDD VSS sg13g2_FILL8
XSTDFILL81_1456 VDD VSS sg13g2_FILL8
XSTDFILL81_1464 VDD VSS sg13g2_FILL8
XSTDFILL81_1472 VDD VSS sg13g2_FILL8
XSTDFILL81_1480 VDD VSS sg13g2_FILL8
XSTDFILL81_1488 VDD VSS sg13g2_FILL8
XSTDFILL81_1496 VDD VSS sg13g2_FILL8
XSTDFILL81_1504 VDD VSS sg13g2_FILL8
XSTDFILL81_1512 VDD VSS sg13g2_FILL8
XSTDFILL81_1520 VDD VSS sg13g2_FILL8
XSTDFILL81_1528 VDD VSS sg13g2_FILL2
XSTDFILL81_1530 VDD VSS sg13g2_FILL1
XSTDFILL82_0 VDD VSS sg13g2_FILL8
XSTDFILL82_8 VDD VSS sg13g2_FILL8
XSTDFILL82_16 VDD VSS sg13g2_FILL8
XSTDFILL82_24 VDD VSS sg13g2_FILL8
XSTDFILL82_32 VDD VSS sg13g2_FILL8
XSTDFILL82_40 VDD VSS sg13g2_FILL8
XSTDFILL82_48 VDD VSS sg13g2_FILL8
XSTDFILL82_56 VDD VSS sg13g2_FILL8
XSTDFILL82_64 VDD VSS sg13g2_FILL8
XSTDFILL82_72 VDD VSS sg13g2_FILL8
XSTDFILL82_80 VDD VSS sg13g2_FILL8
XSTDFILL82_88 VDD VSS sg13g2_FILL8
XSTDFILL82_96 VDD VSS sg13g2_FILL8
XSTDFILL82_104 VDD VSS sg13g2_FILL8
XSTDFILL82_112 VDD VSS sg13g2_FILL8
XSTDFILL82_120 VDD VSS sg13g2_FILL8
XSTDFILL82_128 VDD VSS sg13g2_FILL8
XSTDFILL82_136 VDD VSS sg13g2_FILL8
XSTDFILL82_144 VDD VSS sg13g2_FILL8
XSTDFILL82_152 VDD VSS sg13g2_FILL8
XSTDFILL82_160 VDD VSS sg13g2_FILL8
XSTDFILL82_168 VDD VSS sg13g2_FILL8
XSTDFILL82_176 VDD VSS sg13g2_FILL8
XSTDFILL82_184 VDD VSS sg13g2_FILL8
XSTDFILL82_192 VDD VSS sg13g2_FILL8
XSTDFILL82_200 VDD VSS sg13g2_FILL8
XSTDFILL82_208 VDD VSS sg13g2_FILL8
XSTDFILL82_216 VDD VSS sg13g2_FILL8
XSTDFILL82_224 VDD VSS sg13g2_FILL8
XSTDFILL82_232 VDD VSS sg13g2_FILL8
XSTDFILL82_240 VDD VSS sg13g2_FILL8
XSTDFILL82_248 VDD VSS sg13g2_FILL8
XSTDFILL82_256 VDD VSS sg13g2_FILL8
XSTDFILL82_264 VDD VSS sg13g2_FILL8
XSTDFILL82_272 VDD VSS sg13g2_FILL8
XSTDFILL82_280 VDD VSS sg13g2_FILL8
XSTDFILL82_288 VDD VSS sg13g2_FILL8
XSTDFILL82_296 VDD VSS sg13g2_FILL8
XSTDFILL82_304 VDD VSS sg13g2_FILL8
XSTDFILL82_312 VDD VSS sg13g2_FILL8
XSTDFILL82_320 VDD VSS sg13g2_FILL8
XSTDFILL82_328 VDD VSS sg13g2_FILL8
XSTDFILL82_336 VDD VSS sg13g2_FILL8
XSTDFILL82_344 VDD VSS sg13g2_FILL8
XSTDFILL82_352 VDD VSS sg13g2_FILL8
XSTDFILL82_360 VDD VSS sg13g2_FILL8
XSTDFILL82_368 VDD VSS sg13g2_FILL8
XSTDFILL82_376 VDD VSS sg13g2_FILL8
XSTDFILL82_384 VDD VSS sg13g2_FILL8
XSTDFILL82_392 VDD VSS sg13g2_FILL8
XSTDFILL82_400 VDD VSS sg13g2_FILL8
XSTDFILL82_408 VDD VSS sg13g2_FILL8
XSTDFILL82_416 VDD VSS sg13g2_FILL8
XSTDFILL82_424 VDD VSS sg13g2_FILL8
XSTDFILL82_432 VDD VSS sg13g2_FILL8
XSTDFILL82_440 VDD VSS sg13g2_FILL8
XSTDFILL82_448 VDD VSS sg13g2_FILL8
XSTDFILL82_456 VDD VSS sg13g2_FILL8
XSTDFILL82_464 VDD VSS sg13g2_FILL8
XSTDFILL82_472 VDD VSS sg13g2_FILL8
XSTDFILL82_480 VDD VSS sg13g2_FILL8
XSTDFILL82_488 VDD VSS sg13g2_FILL8
XSTDFILL82_496 VDD VSS sg13g2_FILL8
XSTDFILL82_504 VDD VSS sg13g2_FILL8
XSTDFILL82_512 VDD VSS sg13g2_FILL8
XSTDFILL82_520 VDD VSS sg13g2_FILL8
XSTDFILL82_528 VDD VSS sg13g2_FILL8
XSTDFILL82_536 VDD VSS sg13g2_FILL8
XSTDFILL82_544 VDD VSS sg13g2_FILL8
XSTDFILL82_552 VDD VSS sg13g2_FILL8
XSTDFILL82_560 VDD VSS sg13g2_FILL8
XSTDFILL82_568 VDD VSS sg13g2_FILL8
XSTDFILL82_576 VDD VSS sg13g2_FILL8
XSTDFILL82_584 VDD VSS sg13g2_FILL8
XSTDFILL82_592 VDD VSS sg13g2_FILL8
XSTDFILL82_600 VDD VSS sg13g2_FILL8
XSTDFILL82_608 VDD VSS sg13g2_FILL8
XSTDFILL82_616 VDD VSS sg13g2_FILL8
XSTDFILL82_624 VDD VSS sg13g2_FILL8
XSTDFILL82_632 VDD VSS sg13g2_FILL8
XSTDFILL82_640 VDD VSS sg13g2_FILL8
XSTDFILL82_648 VDD VSS sg13g2_FILL8
XSTDFILL82_656 VDD VSS sg13g2_FILL8
XSTDFILL82_664 VDD VSS sg13g2_FILL8
XSTDFILL82_672 VDD VSS sg13g2_FILL8
XSTDFILL82_680 VDD VSS sg13g2_FILL8
XSTDFILL82_688 VDD VSS sg13g2_FILL8
XSTDFILL82_696 VDD VSS sg13g2_FILL8
XSTDFILL82_704 VDD VSS sg13g2_FILL8
XSTDFILL82_712 VDD VSS sg13g2_FILL8
XSTDFILL82_720 VDD VSS sg13g2_FILL8
XSTDFILL82_728 VDD VSS sg13g2_FILL8
XSTDFILL82_736 VDD VSS sg13g2_FILL8
XSTDFILL82_744 VDD VSS sg13g2_FILL8
XSTDFILL82_752 VDD VSS sg13g2_FILL8
XSTDFILL82_760 VDD VSS sg13g2_FILL8
XSTDFILL82_768 VDD VSS sg13g2_FILL8
XSTDFILL82_776 VDD VSS sg13g2_FILL8
XSTDFILL82_784 VDD VSS sg13g2_FILL8
XSTDFILL82_792 VDD VSS sg13g2_FILL8
XSTDFILL82_800 VDD VSS sg13g2_FILL8
XSTDFILL82_808 VDD VSS sg13g2_FILL8
XSTDFILL82_816 VDD VSS sg13g2_FILL8
XSTDFILL82_824 VDD VSS sg13g2_FILL8
XSTDFILL82_832 VDD VSS sg13g2_FILL8
XSTDFILL82_840 VDD VSS sg13g2_FILL8
XSTDFILL82_848 VDD VSS sg13g2_FILL8
XSTDFILL82_856 VDD VSS sg13g2_FILL8
XSTDFILL82_864 VDD VSS sg13g2_FILL8
XSTDFILL82_872 VDD VSS sg13g2_FILL8
XSTDFILL82_880 VDD VSS sg13g2_FILL8
XSTDFILL82_888 VDD VSS sg13g2_FILL8
XSTDFILL82_896 VDD VSS sg13g2_FILL8
XSTDFILL82_904 VDD VSS sg13g2_FILL8
XSTDFILL82_912 VDD VSS sg13g2_FILL8
XSTDFILL82_920 VDD VSS sg13g2_FILL8
XSTDFILL82_928 VDD VSS sg13g2_FILL8
XSTDFILL82_936 VDD VSS sg13g2_FILL8
XSTDFILL82_944 VDD VSS sg13g2_FILL8
XSTDFILL82_952 VDD VSS sg13g2_FILL8
XSTDFILL82_960 VDD VSS sg13g2_FILL8
XSTDFILL82_968 VDD VSS sg13g2_FILL8
XSTDFILL82_976 VDD VSS sg13g2_FILL8
XSTDFILL82_984 VDD VSS sg13g2_FILL8
XSTDFILL82_992 VDD VSS sg13g2_FILL8
XSTDFILL82_1000 VDD VSS sg13g2_FILL8
XSTDFILL82_1008 VDD VSS sg13g2_FILL8
XSTDFILL82_1016 VDD VSS sg13g2_FILL8
XSTDFILL82_1024 VDD VSS sg13g2_FILL8
XSTDFILL82_1032 VDD VSS sg13g2_FILL8
XSTDFILL82_1040 VDD VSS sg13g2_FILL8
XSTDFILL82_1048 VDD VSS sg13g2_FILL8
XSTDFILL82_1056 VDD VSS sg13g2_FILL8
XSTDFILL82_1064 VDD VSS sg13g2_FILL8
XSTDFILL82_1072 VDD VSS sg13g2_FILL8
XSTDFILL82_1080 VDD VSS sg13g2_FILL8
XSTDFILL82_1088 VDD VSS sg13g2_FILL8
XSTDFILL82_1096 VDD VSS sg13g2_FILL8
XSTDFILL82_1104 VDD VSS sg13g2_FILL8
XSTDFILL82_1112 VDD VSS sg13g2_FILL8
XSTDFILL82_1120 VDD VSS sg13g2_FILL8
XSTDFILL82_1128 VDD VSS sg13g2_FILL8
XSTDFILL82_1136 VDD VSS sg13g2_FILL8
XSTDFILL82_1144 VDD VSS sg13g2_FILL8
XSTDFILL82_1152 VDD VSS sg13g2_FILL8
XSTDFILL82_1160 VDD VSS sg13g2_FILL8
XSTDFILL82_1168 VDD VSS sg13g2_FILL8
XSTDFILL82_1176 VDD VSS sg13g2_FILL8
XSTDFILL82_1184 VDD VSS sg13g2_FILL8
XSTDFILL82_1192 VDD VSS sg13g2_FILL8
XSTDFILL82_1200 VDD VSS sg13g2_FILL8
XSTDFILL82_1208 VDD VSS sg13g2_FILL8
XSTDFILL82_1216 VDD VSS sg13g2_FILL8
XSTDFILL82_1224 VDD VSS sg13g2_FILL8
XSTDFILL82_1232 VDD VSS sg13g2_FILL8
XSTDFILL82_1240 VDD VSS sg13g2_FILL8
XSTDFILL82_1248 VDD VSS sg13g2_FILL8
XSTDFILL82_1256 VDD VSS sg13g2_FILL8
XSTDFILL82_1264 VDD VSS sg13g2_FILL8
XSTDFILL82_1272 VDD VSS sg13g2_FILL8
XSTDFILL82_1280 VDD VSS sg13g2_FILL8
XSTDFILL82_1288 VDD VSS sg13g2_FILL8
XSTDFILL82_1296 VDD VSS sg13g2_FILL8
XSTDFILL82_1304 VDD VSS sg13g2_FILL8
XSTDFILL82_1312 VDD VSS sg13g2_FILL8
XSTDFILL82_1320 VDD VSS sg13g2_FILL8
XSTDFILL82_1328 VDD VSS sg13g2_FILL8
XSTDFILL82_1336 VDD VSS sg13g2_FILL8
XSTDFILL82_1344 VDD VSS sg13g2_FILL8
XSTDFILL82_1352 VDD VSS sg13g2_FILL8
XSTDFILL82_1360 VDD VSS sg13g2_FILL8
XSTDFILL82_1368 VDD VSS sg13g2_FILL8
XSTDFILL82_1376 VDD VSS sg13g2_FILL8
XSTDFILL82_1384 VDD VSS sg13g2_FILL8
XSTDFILL82_1392 VDD VSS sg13g2_FILL8
XSTDFILL82_1400 VDD VSS sg13g2_FILL8
XSTDFILL82_1408 VDD VSS sg13g2_FILL8
XSTDFILL82_1416 VDD VSS sg13g2_FILL8
XSTDFILL82_1424 VDD VSS sg13g2_FILL8
XSTDFILL82_1432 VDD VSS sg13g2_FILL8
XSTDFILL82_1440 VDD VSS sg13g2_FILL8
XSTDFILL82_1448 VDD VSS sg13g2_FILL8
XSTDFILL82_1456 VDD VSS sg13g2_FILL8
XSTDFILL82_1464 VDD VSS sg13g2_FILL8
XSTDFILL82_1472 VDD VSS sg13g2_FILL8
XSTDFILL82_1480 VDD VSS sg13g2_FILL8
XSTDFILL82_1488 VDD VSS sg13g2_FILL8
XSTDFILL82_1496 VDD VSS sg13g2_FILL8
XSTDFILL82_1504 VDD VSS sg13g2_FILL8
XSTDFILL82_1512 VDD VSS sg13g2_FILL8
XSTDFILL82_1520 VDD VSS sg13g2_FILL8
XSTDFILL82_1528 VDD VSS sg13g2_FILL2
XSTDFILL82_1530 VDD VSS sg13g2_FILL1
XSTDFILL83_0 VDD VSS sg13g2_FILL8
XSTDFILL83_8 VDD VSS sg13g2_FILL8
XSTDFILL83_16 VDD VSS sg13g2_FILL8
XSTDFILL83_24 VDD VSS sg13g2_FILL8
XSTDFILL83_32 VDD VSS sg13g2_FILL8
XSTDFILL83_40 VDD VSS sg13g2_FILL8
XSTDFILL83_48 VDD VSS sg13g2_FILL8
XSTDFILL83_56 VDD VSS sg13g2_FILL8
XSTDFILL83_64 VDD VSS sg13g2_FILL8
XSTDFILL83_72 VDD VSS sg13g2_FILL8
XSTDFILL83_80 VDD VSS sg13g2_FILL8
XSTDFILL83_88 VDD VSS sg13g2_FILL8
XSTDFILL83_96 VDD VSS sg13g2_FILL8
XSTDFILL83_104 VDD VSS sg13g2_FILL8
XSTDFILL83_112 VDD VSS sg13g2_FILL8
XSTDFILL83_120 VDD VSS sg13g2_FILL8
XSTDFILL83_128 VDD VSS sg13g2_FILL8
XSTDFILL83_136 VDD VSS sg13g2_FILL8
XSTDFILL83_144 VDD VSS sg13g2_FILL8
XSTDFILL83_152 VDD VSS sg13g2_FILL8
XSTDFILL83_160 VDD VSS sg13g2_FILL8
XSTDFILL83_168 VDD VSS sg13g2_FILL8
XSTDFILL83_176 VDD VSS sg13g2_FILL8
XSTDFILL83_184 VDD VSS sg13g2_FILL8
XSTDFILL83_192 VDD VSS sg13g2_FILL8
XSTDFILL83_200 VDD VSS sg13g2_FILL8
XSTDFILL83_208 VDD VSS sg13g2_FILL8
XSTDFILL83_216 VDD VSS sg13g2_FILL8
XSTDFILL83_224 VDD VSS sg13g2_FILL8
XSTDFILL83_232 VDD VSS sg13g2_FILL8
XSTDFILL83_240 VDD VSS sg13g2_FILL8
XSTDFILL83_248 VDD VSS sg13g2_FILL8
XSTDFILL83_256 VDD VSS sg13g2_FILL8
XSTDFILL83_264 VDD VSS sg13g2_FILL8
XSTDFILL83_272 VDD VSS sg13g2_FILL8
XSTDFILL83_280 VDD VSS sg13g2_FILL8
XSTDFILL83_288 VDD VSS sg13g2_FILL8
XSTDFILL83_296 VDD VSS sg13g2_FILL8
XSTDFILL83_304 VDD VSS sg13g2_FILL8
XSTDFILL83_312 VDD VSS sg13g2_FILL8
XSTDFILL83_320 VDD VSS sg13g2_FILL8
XSTDFILL83_328 VDD VSS sg13g2_FILL8
XSTDFILL83_336 VDD VSS sg13g2_FILL8
XSTDFILL83_344 VDD VSS sg13g2_FILL8
XSTDFILL83_352 VDD VSS sg13g2_FILL8
XSTDFILL83_360 VDD VSS sg13g2_FILL8
XSTDFILL83_368 VDD VSS sg13g2_FILL8
XSTDFILL83_376 VDD VSS sg13g2_FILL8
XSTDFILL83_384 VDD VSS sg13g2_FILL8
XSTDFILL83_392 VDD VSS sg13g2_FILL8
XSTDFILL83_400 VDD VSS sg13g2_FILL8
XSTDFILL83_408 VDD VSS sg13g2_FILL8
XSTDFILL83_416 VDD VSS sg13g2_FILL8
XSTDFILL83_424 VDD VSS sg13g2_FILL8
XSTDFILL83_432 VDD VSS sg13g2_FILL8
XSTDFILL83_440 VDD VSS sg13g2_FILL8
XSTDFILL83_448 VDD VSS sg13g2_FILL8
XSTDFILL83_456 VDD VSS sg13g2_FILL8
XSTDFILL83_464 VDD VSS sg13g2_FILL8
XSTDFILL83_472 VDD VSS sg13g2_FILL8
XSTDFILL83_480 VDD VSS sg13g2_FILL8
XSTDFILL83_488 VDD VSS sg13g2_FILL8
XSTDFILL83_496 VDD VSS sg13g2_FILL8
XSTDFILL83_504 VDD VSS sg13g2_FILL8
XSTDFILL83_512 VDD VSS sg13g2_FILL8
XSTDFILL83_520 VDD VSS sg13g2_FILL8
XSTDFILL83_528 VDD VSS sg13g2_FILL8
XSTDFILL83_536 VDD VSS sg13g2_FILL8
XSTDFILL83_544 VDD VSS sg13g2_FILL8
XSTDFILL83_552 VDD VSS sg13g2_FILL8
XSTDFILL83_560 VDD VSS sg13g2_FILL8
XSTDFILL83_568 VDD VSS sg13g2_FILL8
XSTDFILL83_576 VDD VSS sg13g2_FILL8
XSTDFILL83_584 VDD VSS sg13g2_FILL8
XSTDFILL83_592 VDD VSS sg13g2_FILL8
XSTDFILL83_600 VDD VSS sg13g2_FILL8
XSTDFILL83_608 VDD VSS sg13g2_FILL8
XSTDFILL83_616 VDD VSS sg13g2_FILL8
XSTDFILL83_624 VDD VSS sg13g2_FILL8
XSTDFILL83_632 VDD VSS sg13g2_FILL8
XSTDFILL83_640 VDD VSS sg13g2_FILL8
XSTDFILL83_648 VDD VSS sg13g2_FILL8
XSTDFILL83_656 VDD VSS sg13g2_FILL8
XSTDFILL83_664 VDD VSS sg13g2_FILL8
XSTDFILL83_672 VDD VSS sg13g2_FILL8
XSTDFILL83_680 VDD VSS sg13g2_FILL8
XSTDFILL83_688 VDD VSS sg13g2_FILL8
XSTDFILL83_696 VDD VSS sg13g2_FILL8
XSTDFILL83_704 VDD VSS sg13g2_FILL8
XSTDFILL83_712 VDD VSS sg13g2_FILL8
XSTDFILL83_720 VDD VSS sg13g2_FILL8
XSTDFILL83_728 VDD VSS sg13g2_FILL8
XSTDFILL83_736 VDD VSS sg13g2_FILL8
XSTDFILL83_744 VDD VSS sg13g2_FILL8
XSTDFILL83_752 VDD VSS sg13g2_FILL8
XSTDFILL83_760 VDD VSS sg13g2_FILL8
XSTDFILL83_768 VDD VSS sg13g2_FILL8
XSTDFILL83_776 VDD VSS sg13g2_FILL8
XSTDFILL83_784 VDD VSS sg13g2_FILL8
XSTDFILL83_792 VDD VSS sg13g2_FILL8
XSTDFILL83_800 VDD VSS sg13g2_FILL8
XSTDFILL83_808 VDD VSS sg13g2_FILL8
XSTDFILL83_816 VDD VSS sg13g2_FILL8
XSTDFILL83_824 VDD VSS sg13g2_FILL8
XSTDFILL83_832 VDD VSS sg13g2_FILL8
XSTDFILL83_840 VDD VSS sg13g2_FILL8
XSTDFILL83_848 VDD VSS sg13g2_FILL8
XSTDFILL83_856 VDD VSS sg13g2_FILL8
XSTDFILL83_864 VDD VSS sg13g2_FILL8
XSTDFILL83_872 VDD VSS sg13g2_FILL8
XSTDFILL83_880 VDD VSS sg13g2_FILL8
XSTDFILL83_888 VDD VSS sg13g2_FILL8
XSTDFILL83_896 VDD VSS sg13g2_FILL8
XSTDFILL83_904 VDD VSS sg13g2_FILL8
XSTDFILL83_912 VDD VSS sg13g2_FILL8
XSTDFILL83_920 VDD VSS sg13g2_FILL8
XSTDFILL83_928 VDD VSS sg13g2_FILL8
XSTDFILL83_936 VDD VSS sg13g2_FILL8
XSTDFILL83_944 VDD VSS sg13g2_FILL8
XSTDFILL83_952 VDD VSS sg13g2_FILL8
XSTDFILL83_960 VDD VSS sg13g2_FILL8
XSTDFILL83_968 VDD VSS sg13g2_FILL8
XSTDFILL83_976 VDD VSS sg13g2_FILL8
XSTDFILL83_984 VDD VSS sg13g2_FILL8
XSTDFILL83_992 VDD VSS sg13g2_FILL8
XSTDFILL83_1000 VDD VSS sg13g2_FILL8
XSTDFILL83_1008 VDD VSS sg13g2_FILL8
XSTDFILL83_1016 VDD VSS sg13g2_FILL8
XSTDFILL83_1024 VDD VSS sg13g2_FILL8
XSTDFILL83_1032 VDD VSS sg13g2_FILL8
XSTDFILL83_1040 VDD VSS sg13g2_FILL8
XSTDFILL83_1048 VDD VSS sg13g2_FILL8
XSTDFILL83_1056 VDD VSS sg13g2_FILL8
XSTDFILL83_1064 VDD VSS sg13g2_FILL8
XSTDFILL83_1072 VDD VSS sg13g2_FILL8
XSTDFILL83_1080 VDD VSS sg13g2_FILL8
XSTDFILL83_1088 VDD VSS sg13g2_FILL8
XSTDFILL83_1096 VDD VSS sg13g2_FILL8
XSTDFILL83_1104 VDD VSS sg13g2_FILL8
XSTDFILL83_1112 VDD VSS sg13g2_FILL8
XSTDFILL83_1120 VDD VSS sg13g2_FILL8
XSTDFILL83_1128 VDD VSS sg13g2_FILL8
XSTDFILL83_1136 VDD VSS sg13g2_FILL8
XSTDFILL83_1144 VDD VSS sg13g2_FILL8
XSTDFILL83_1152 VDD VSS sg13g2_FILL8
XSTDFILL83_1160 VDD VSS sg13g2_FILL8
XSTDFILL83_1168 VDD VSS sg13g2_FILL8
XSTDFILL83_1176 VDD VSS sg13g2_FILL8
XSTDFILL83_1184 VDD VSS sg13g2_FILL8
XSTDFILL83_1192 VDD VSS sg13g2_FILL8
XSTDFILL83_1200 VDD VSS sg13g2_FILL8
XSTDFILL83_1208 VDD VSS sg13g2_FILL8
XSTDFILL83_1216 VDD VSS sg13g2_FILL8
XSTDFILL83_1224 VDD VSS sg13g2_FILL8
XSTDFILL83_1232 VDD VSS sg13g2_FILL8
XSTDFILL83_1240 VDD VSS sg13g2_FILL8
XSTDFILL83_1248 VDD VSS sg13g2_FILL8
XSTDFILL83_1256 VDD VSS sg13g2_FILL8
XSTDFILL83_1264 VDD VSS sg13g2_FILL8
XSTDFILL83_1272 VDD VSS sg13g2_FILL8
XSTDFILL83_1280 VDD VSS sg13g2_FILL8
XSTDFILL83_1288 VDD VSS sg13g2_FILL8
XSTDFILL83_1296 VDD VSS sg13g2_FILL8
XSTDFILL83_1304 VDD VSS sg13g2_FILL8
XSTDFILL83_1312 VDD VSS sg13g2_FILL8
XSTDFILL83_1320 VDD VSS sg13g2_FILL8
XSTDFILL83_1328 VDD VSS sg13g2_FILL8
XSTDFILL83_1336 VDD VSS sg13g2_FILL8
XSTDFILL83_1344 VDD VSS sg13g2_FILL8
XSTDFILL83_1352 VDD VSS sg13g2_FILL8
XSTDFILL83_1360 VDD VSS sg13g2_FILL8
XSTDFILL83_1368 VDD VSS sg13g2_FILL8
XSTDFILL83_1376 VDD VSS sg13g2_FILL8
XSTDFILL83_1384 VDD VSS sg13g2_FILL8
XSTDFILL83_1392 VDD VSS sg13g2_FILL8
XSTDFILL83_1400 VDD VSS sg13g2_FILL8
XSTDFILL83_1408 VDD VSS sg13g2_FILL8
XSTDFILL83_1416 VDD VSS sg13g2_FILL8
XSTDFILL83_1424 VDD VSS sg13g2_FILL8
XSTDFILL83_1432 VDD VSS sg13g2_FILL8
XSTDFILL83_1440 VDD VSS sg13g2_FILL8
XSTDFILL83_1448 VDD VSS sg13g2_FILL8
XSTDFILL83_1456 VDD VSS sg13g2_FILL8
XSTDFILL83_1464 VDD VSS sg13g2_FILL8
XSTDFILL83_1472 VDD VSS sg13g2_FILL8
XSTDFILL83_1480 VDD VSS sg13g2_FILL8
XSTDFILL83_1488 VDD VSS sg13g2_FILL8
XSTDFILL83_1496 VDD VSS sg13g2_FILL8
XSTDFILL83_1504 VDD VSS sg13g2_FILL8
XSTDFILL83_1512 VDD VSS sg13g2_FILL8
XSTDFILL83_1520 VDD VSS sg13g2_FILL8
XSTDFILL83_1528 VDD VSS sg13g2_FILL2
XSTDFILL83_1530 VDD VSS sg13g2_FILL1
XSTDFILL84_0 VDD VSS sg13g2_FILL8
XSTDFILL84_8 VDD VSS sg13g2_FILL8
XSTDFILL84_16 VDD VSS sg13g2_FILL8
XSTDFILL84_24 VDD VSS sg13g2_FILL8
XSTDFILL84_32 VDD VSS sg13g2_FILL8
XSTDFILL84_40 VDD VSS sg13g2_FILL8
XSTDFILL84_48 VDD VSS sg13g2_FILL8
XSTDFILL84_56 VDD VSS sg13g2_FILL8
XSTDFILL84_64 VDD VSS sg13g2_FILL8
XSTDFILL84_72 VDD VSS sg13g2_FILL8
XSTDFILL84_80 VDD VSS sg13g2_FILL8
XSTDFILL84_88 VDD VSS sg13g2_FILL8
XSTDFILL84_96 VDD VSS sg13g2_FILL8
XSTDFILL84_104 VDD VSS sg13g2_FILL8
XSTDFILL84_112 VDD VSS sg13g2_FILL8
XSTDFILL84_120 VDD VSS sg13g2_FILL8
XSTDFILL84_128 VDD VSS sg13g2_FILL8
XSTDFILL84_136 VDD VSS sg13g2_FILL8
XSTDFILL84_144 VDD VSS sg13g2_FILL8
XSTDFILL84_152 VDD VSS sg13g2_FILL8
XSTDFILL84_160 VDD VSS sg13g2_FILL8
XSTDFILL84_168 VDD VSS sg13g2_FILL8
XSTDFILL84_176 VDD VSS sg13g2_FILL8
XSTDFILL84_184 VDD VSS sg13g2_FILL8
XSTDFILL84_192 VDD VSS sg13g2_FILL8
XSTDFILL84_200 VDD VSS sg13g2_FILL8
XSTDFILL84_208 VDD VSS sg13g2_FILL8
XSTDFILL84_216 VDD VSS sg13g2_FILL8
XSTDFILL84_224 VDD VSS sg13g2_FILL8
XSTDFILL84_232 VDD VSS sg13g2_FILL8
XSTDFILL84_240 VDD VSS sg13g2_FILL8
XSTDFILL84_248 VDD VSS sg13g2_FILL8
XSTDFILL84_256 VDD VSS sg13g2_FILL8
XSTDFILL84_264 VDD VSS sg13g2_FILL8
XSTDFILL84_272 VDD VSS sg13g2_FILL8
XSTDFILL84_280 VDD VSS sg13g2_FILL8
XSTDFILL84_288 VDD VSS sg13g2_FILL8
XSTDFILL84_296 VDD VSS sg13g2_FILL8
XSTDFILL84_304 VDD VSS sg13g2_FILL8
XSTDFILL84_312 VDD VSS sg13g2_FILL8
XSTDFILL84_320 VDD VSS sg13g2_FILL8
XSTDFILL84_328 VDD VSS sg13g2_FILL8
XSTDFILL84_336 VDD VSS sg13g2_FILL8
XSTDFILL84_344 VDD VSS sg13g2_FILL8
XSTDFILL84_352 VDD VSS sg13g2_FILL8
XSTDFILL84_360 VDD VSS sg13g2_FILL8
XSTDFILL84_368 VDD VSS sg13g2_FILL8
XSTDFILL84_376 VDD VSS sg13g2_FILL8
XSTDFILL84_384 VDD VSS sg13g2_FILL8
XSTDFILL84_392 VDD VSS sg13g2_FILL8
XSTDFILL84_400 VDD VSS sg13g2_FILL8
XSTDFILL84_408 VDD VSS sg13g2_FILL8
XSTDFILL84_416 VDD VSS sg13g2_FILL8
XSTDFILL84_424 VDD VSS sg13g2_FILL8
XSTDFILL84_432 VDD VSS sg13g2_FILL8
XSTDFILL84_440 VDD VSS sg13g2_FILL8
XSTDFILL84_448 VDD VSS sg13g2_FILL8
XSTDFILL84_456 VDD VSS sg13g2_FILL8
XSTDFILL84_464 VDD VSS sg13g2_FILL8
XSTDFILL84_472 VDD VSS sg13g2_FILL8
XSTDFILL84_480 VDD VSS sg13g2_FILL8
XSTDFILL84_488 VDD VSS sg13g2_FILL8
XSTDFILL84_496 VDD VSS sg13g2_FILL8
XSTDFILL84_504 VDD VSS sg13g2_FILL8
XSTDFILL84_512 VDD VSS sg13g2_FILL8
XSTDFILL84_520 VDD VSS sg13g2_FILL8
XSTDFILL84_528 VDD VSS sg13g2_FILL8
XSTDFILL84_536 VDD VSS sg13g2_FILL8
XSTDFILL84_544 VDD VSS sg13g2_FILL8
XSTDFILL84_552 VDD VSS sg13g2_FILL8
XSTDFILL84_560 VDD VSS sg13g2_FILL8
XSTDFILL84_568 VDD VSS sg13g2_FILL8
XSTDFILL84_576 VDD VSS sg13g2_FILL8
XSTDFILL84_584 VDD VSS sg13g2_FILL8
XSTDFILL84_592 VDD VSS sg13g2_FILL8
XSTDFILL84_600 VDD VSS sg13g2_FILL8
XSTDFILL84_608 VDD VSS sg13g2_FILL8
XSTDFILL84_616 VDD VSS sg13g2_FILL8
XSTDFILL84_624 VDD VSS sg13g2_FILL8
XSTDFILL84_632 VDD VSS sg13g2_FILL8
XSTDFILL84_640 VDD VSS sg13g2_FILL8
XSTDFILL84_648 VDD VSS sg13g2_FILL8
XSTDFILL84_656 VDD VSS sg13g2_FILL8
XSTDFILL84_664 VDD VSS sg13g2_FILL8
XSTDFILL84_672 VDD VSS sg13g2_FILL8
XSTDFILL84_680 VDD VSS sg13g2_FILL8
XSTDFILL84_688 VDD VSS sg13g2_FILL8
XSTDFILL84_696 VDD VSS sg13g2_FILL8
XSTDFILL84_704 VDD VSS sg13g2_FILL8
XSTDFILL84_712 VDD VSS sg13g2_FILL8
XSTDFILL84_720 VDD VSS sg13g2_FILL8
XSTDFILL84_728 VDD VSS sg13g2_FILL8
XSTDFILL84_736 VDD VSS sg13g2_FILL8
XSTDFILL84_744 VDD VSS sg13g2_FILL8
XSTDFILL84_752 VDD VSS sg13g2_FILL8
XSTDFILL84_760 VDD VSS sg13g2_FILL8
XSTDFILL84_768 VDD VSS sg13g2_FILL8
XSTDFILL84_776 VDD VSS sg13g2_FILL8
XSTDFILL84_784 VDD VSS sg13g2_FILL8
XSTDFILL84_792 VDD VSS sg13g2_FILL8
XSTDFILL84_800 VDD VSS sg13g2_FILL8
XSTDFILL84_808 VDD VSS sg13g2_FILL8
XSTDFILL84_816 VDD VSS sg13g2_FILL8
XSTDFILL84_824 VDD VSS sg13g2_FILL8
XSTDFILL84_832 VDD VSS sg13g2_FILL8
XSTDFILL84_840 VDD VSS sg13g2_FILL8
XSTDFILL84_848 VDD VSS sg13g2_FILL8
XSTDFILL84_856 VDD VSS sg13g2_FILL8
XSTDFILL84_864 VDD VSS sg13g2_FILL8
XSTDFILL84_872 VDD VSS sg13g2_FILL8
XSTDFILL84_880 VDD VSS sg13g2_FILL8
XSTDFILL84_888 VDD VSS sg13g2_FILL8
XSTDFILL84_896 VDD VSS sg13g2_FILL8
XSTDFILL84_904 VDD VSS sg13g2_FILL8
XSTDFILL84_912 VDD VSS sg13g2_FILL8
XSTDFILL84_920 VDD VSS sg13g2_FILL8
XSTDFILL84_928 VDD VSS sg13g2_FILL8
XSTDFILL84_936 VDD VSS sg13g2_FILL8
XSTDFILL84_944 VDD VSS sg13g2_FILL8
XSTDFILL84_952 VDD VSS sg13g2_FILL8
XSTDFILL84_960 VDD VSS sg13g2_FILL8
XSTDFILL84_968 VDD VSS sg13g2_FILL8
XSTDFILL84_976 VDD VSS sg13g2_FILL8
XSTDFILL84_984 VDD VSS sg13g2_FILL8
XSTDFILL84_992 VDD VSS sg13g2_FILL8
XSTDFILL84_1000 VDD VSS sg13g2_FILL8
XSTDFILL84_1008 VDD VSS sg13g2_FILL8
XSTDFILL84_1016 VDD VSS sg13g2_FILL8
XSTDFILL84_1024 VDD VSS sg13g2_FILL8
XSTDFILL84_1032 VDD VSS sg13g2_FILL8
XSTDFILL84_1040 VDD VSS sg13g2_FILL8
XSTDFILL84_1048 VDD VSS sg13g2_FILL8
XSTDFILL84_1056 VDD VSS sg13g2_FILL8
XSTDFILL84_1064 VDD VSS sg13g2_FILL8
XSTDFILL84_1072 VDD VSS sg13g2_FILL8
XSTDFILL84_1080 VDD VSS sg13g2_FILL8
XSTDFILL84_1088 VDD VSS sg13g2_FILL8
XSTDFILL84_1096 VDD VSS sg13g2_FILL8
XSTDFILL84_1104 VDD VSS sg13g2_FILL8
XSTDFILL84_1112 VDD VSS sg13g2_FILL8
XSTDFILL84_1120 VDD VSS sg13g2_FILL8
XSTDFILL84_1128 VDD VSS sg13g2_FILL8
XSTDFILL84_1136 VDD VSS sg13g2_FILL8
XSTDFILL84_1144 VDD VSS sg13g2_FILL8
XSTDFILL84_1152 VDD VSS sg13g2_FILL8
XSTDFILL84_1160 VDD VSS sg13g2_FILL8
XSTDFILL84_1168 VDD VSS sg13g2_FILL8
XSTDFILL84_1176 VDD VSS sg13g2_FILL8
XSTDFILL84_1184 VDD VSS sg13g2_FILL8
XSTDFILL84_1192 VDD VSS sg13g2_FILL8
XSTDFILL84_1200 VDD VSS sg13g2_FILL8
XSTDFILL84_1208 VDD VSS sg13g2_FILL8
XSTDFILL84_1216 VDD VSS sg13g2_FILL8
XSTDFILL84_1224 VDD VSS sg13g2_FILL8
XSTDFILL84_1232 VDD VSS sg13g2_FILL8
XSTDFILL84_1240 VDD VSS sg13g2_FILL8
XSTDFILL84_1248 VDD VSS sg13g2_FILL8
XSTDFILL84_1256 VDD VSS sg13g2_FILL8
XSTDFILL84_1264 VDD VSS sg13g2_FILL8
XSTDFILL84_1272 VDD VSS sg13g2_FILL8
XSTDFILL84_1280 VDD VSS sg13g2_FILL8
XSTDFILL84_1288 VDD VSS sg13g2_FILL8
XSTDFILL84_1296 VDD VSS sg13g2_FILL8
XSTDFILL84_1304 VDD VSS sg13g2_FILL8
XSTDFILL84_1312 VDD VSS sg13g2_FILL8
XSTDFILL84_1320 VDD VSS sg13g2_FILL8
XSTDFILL84_1328 VDD VSS sg13g2_FILL8
XSTDFILL84_1336 VDD VSS sg13g2_FILL8
XSTDFILL84_1344 VDD VSS sg13g2_FILL8
XSTDFILL84_1352 VDD VSS sg13g2_FILL8
XSTDFILL84_1360 VDD VSS sg13g2_FILL8
XSTDFILL84_1368 VDD VSS sg13g2_FILL8
XSTDFILL84_1376 VDD VSS sg13g2_FILL8
XSTDFILL84_1384 VDD VSS sg13g2_FILL8
XSTDFILL84_1392 VDD VSS sg13g2_FILL8
XSTDFILL84_1400 VDD VSS sg13g2_FILL8
XSTDFILL84_1408 VDD VSS sg13g2_FILL8
XSTDFILL84_1416 VDD VSS sg13g2_FILL8
XSTDFILL84_1424 VDD VSS sg13g2_FILL8
XSTDFILL84_1432 VDD VSS sg13g2_FILL8
XSTDFILL84_1440 VDD VSS sg13g2_FILL8
XSTDFILL84_1448 VDD VSS sg13g2_FILL8
XSTDFILL84_1456 VDD VSS sg13g2_FILL8
XSTDFILL84_1464 VDD VSS sg13g2_FILL8
XSTDFILL84_1472 VDD VSS sg13g2_FILL8
XSTDFILL84_1480 VDD VSS sg13g2_FILL8
XSTDFILL84_1488 VDD VSS sg13g2_FILL8
XSTDFILL84_1496 VDD VSS sg13g2_FILL8
XSTDFILL84_1504 VDD VSS sg13g2_FILL8
XSTDFILL84_1512 VDD VSS sg13g2_FILL8
XSTDFILL84_1520 VDD VSS sg13g2_FILL8
XSTDFILL84_1528 VDD VSS sg13g2_FILL2
XSTDFILL84_1530 VDD VSS sg13g2_FILL1
XSTDFILL85_0 VDD VSS sg13g2_FILL8
XSTDFILL85_8 VDD VSS sg13g2_FILL8
XSTDFILL85_16 VDD VSS sg13g2_FILL8
XSTDFILL85_24 VDD VSS sg13g2_FILL8
XSTDFILL85_32 VDD VSS sg13g2_FILL8
XSTDFILL85_40 VDD VSS sg13g2_FILL8
XSTDFILL85_48 VDD VSS sg13g2_FILL8
XSTDFILL85_56 VDD VSS sg13g2_FILL8
XSTDFILL85_64 VDD VSS sg13g2_FILL8
XSTDFILL85_72 VDD VSS sg13g2_FILL8
XSTDFILL85_80 VDD VSS sg13g2_FILL8
XSTDFILL85_88 VDD VSS sg13g2_FILL8
XSTDFILL85_96 VDD VSS sg13g2_FILL8
XSTDFILL85_104 VDD VSS sg13g2_FILL8
XSTDFILL85_112 VDD VSS sg13g2_FILL8
XSTDFILL85_120 VDD VSS sg13g2_FILL8
XSTDFILL85_128 VDD VSS sg13g2_FILL8
XSTDFILL85_136 VDD VSS sg13g2_FILL8
XSTDFILL85_144 VDD VSS sg13g2_FILL8
XSTDFILL85_152 VDD VSS sg13g2_FILL8
XSTDFILL85_160 VDD VSS sg13g2_FILL8
XSTDFILL85_168 VDD VSS sg13g2_FILL8
XSTDFILL85_176 VDD VSS sg13g2_FILL8
XSTDFILL85_184 VDD VSS sg13g2_FILL8
XSTDFILL85_192 VDD VSS sg13g2_FILL8
XSTDFILL85_200 VDD VSS sg13g2_FILL8
XSTDFILL85_208 VDD VSS sg13g2_FILL8
XSTDFILL85_216 VDD VSS sg13g2_FILL8
XSTDFILL85_224 VDD VSS sg13g2_FILL8
XSTDFILL85_232 VDD VSS sg13g2_FILL8
XSTDFILL85_240 VDD VSS sg13g2_FILL8
XSTDFILL85_248 VDD VSS sg13g2_FILL8
XSTDFILL85_256 VDD VSS sg13g2_FILL8
XSTDFILL85_264 VDD VSS sg13g2_FILL8
XSTDFILL85_272 VDD VSS sg13g2_FILL8
XSTDFILL85_280 VDD VSS sg13g2_FILL8
XSTDFILL85_288 VDD VSS sg13g2_FILL8
XSTDFILL85_296 VDD VSS sg13g2_FILL8
XSTDFILL85_304 VDD VSS sg13g2_FILL8
XSTDFILL85_312 VDD VSS sg13g2_FILL8
XSTDFILL85_320 VDD VSS sg13g2_FILL8
XSTDFILL85_328 VDD VSS sg13g2_FILL8
XSTDFILL85_336 VDD VSS sg13g2_FILL8
XSTDFILL85_344 VDD VSS sg13g2_FILL8
XSTDFILL85_352 VDD VSS sg13g2_FILL8
XSTDFILL85_360 VDD VSS sg13g2_FILL8
XSTDFILL85_368 VDD VSS sg13g2_FILL8
XSTDFILL85_376 VDD VSS sg13g2_FILL8
XSTDFILL85_384 VDD VSS sg13g2_FILL8
XSTDFILL85_392 VDD VSS sg13g2_FILL8
XSTDFILL85_400 VDD VSS sg13g2_FILL8
XSTDFILL85_408 VDD VSS sg13g2_FILL8
XSTDFILL85_416 VDD VSS sg13g2_FILL8
XSTDFILL85_424 VDD VSS sg13g2_FILL8
XSTDFILL85_432 VDD VSS sg13g2_FILL8
XSTDFILL85_440 VDD VSS sg13g2_FILL8
XSTDFILL85_448 VDD VSS sg13g2_FILL8
XSTDFILL85_456 VDD VSS sg13g2_FILL8
XSTDFILL85_464 VDD VSS sg13g2_FILL8
XSTDFILL85_472 VDD VSS sg13g2_FILL8
XSTDFILL85_480 VDD VSS sg13g2_FILL8
XSTDFILL85_488 VDD VSS sg13g2_FILL8
XSTDFILL85_496 VDD VSS sg13g2_FILL8
XSTDFILL85_504 VDD VSS sg13g2_FILL8
XSTDFILL85_512 VDD VSS sg13g2_FILL8
XSTDFILL85_520 VDD VSS sg13g2_FILL8
XSTDFILL85_528 VDD VSS sg13g2_FILL8
XSTDFILL85_536 VDD VSS sg13g2_FILL8
XSTDFILL85_544 VDD VSS sg13g2_FILL8
XSTDFILL85_552 VDD VSS sg13g2_FILL8
XSTDFILL85_560 VDD VSS sg13g2_FILL8
XSTDFILL85_568 VDD VSS sg13g2_FILL8
XSTDFILL85_576 VDD VSS sg13g2_FILL8
XSTDFILL85_584 VDD VSS sg13g2_FILL8
XSTDFILL85_592 VDD VSS sg13g2_FILL8
XSTDFILL85_600 VDD VSS sg13g2_FILL8
XSTDFILL85_608 VDD VSS sg13g2_FILL8
XSTDFILL85_616 VDD VSS sg13g2_FILL8
XSTDFILL85_624 VDD VSS sg13g2_FILL8
XSTDFILL85_632 VDD VSS sg13g2_FILL8
XSTDFILL85_640 VDD VSS sg13g2_FILL8
XSTDFILL85_648 VDD VSS sg13g2_FILL8
XSTDFILL85_656 VDD VSS sg13g2_FILL8
XSTDFILL85_664 VDD VSS sg13g2_FILL8
XSTDFILL85_672 VDD VSS sg13g2_FILL8
XSTDFILL85_680 VDD VSS sg13g2_FILL8
XSTDFILL85_688 VDD VSS sg13g2_FILL8
XSTDFILL85_696 VDD VSS sg13g2_FILL8
XSTDFILL85_704 VDD VSS sg13g2_FILL8
XSTDFILL85_712 VDD VSS sg13g2_FILL8
XSTDFILL85_720 VDD VSS sg13g2_FILL8
XSTDFILL85_728 VDD VSS sg13g2_FILL8
XSTDFILL85_736 VDD VSS sg13g2_FILL8
XSTDFILL85_744 VDD VSS sg13g2_FILL8
XSTDFILL85_752 VDD VSS sg13g2_FILL8
XSTDFILL85_760 VDD VSS sg13g2_FILL8
XSTDFILL85_768 VDD VSS sg13g2_FILL8
XSTDFILL85_776 VDD VSS sg13g2_FILL8
XSTDFILL85_784 VDD VSS sg13g2_FILL8
XSTDFILL85_792 VDD VSS sg13g2_FILL8
XSTDFILL85_800 VDD VSS sg13g2_FILL8
XSTDFILL85_808 VDD VSS sg13g2_FILL8
XSTDFILL85_816 VDD VSS sg13g2_FILL8
XSTDFILL85_824 VDD VSS sg13g2_FILL8
XSTDFILL85_832 VDD VSS sg13g2_FILL8
XSTDFILL85_840 VDD VSS sg13g2_FILL8
XSTDFILL85_848 VDD VSS sg13g2_FILL8
XSTDFILL85_856 VDD VSS sg13g2_FILL8
XSTDFILL85_864 VDD VSS sg13g2_FILL8
XSTDFILL85_872 VDD VSS sg13g2_FILL8
XSTDFILL85_880 VDD VSS sg13g2_FILL8
XSTDFILL85_888 VDD VSS sg13g2_FILL8
XSTDFILL85_896 VDD VSS sg13g2_FILL8
XSTDFILL85_904 VDD VSS sg13g2_FILL8
XSTDFILL85_912 VDD VSS sg13g2_FILL8
XSTDFILL85_920 VDD VSS sg13g2_FILL8
XSTDFILL85_928 VDD VSS sg13g2_FILL8
XSTDFILL85_936 VDD VSS sg13g2_FILL8
XSTDFILL85_944 VDD VSS sg13g2_FILL8
XSTDFILL85_952 VDD VSS sg13g2_FILL8
XSTDFILL85_960 VDD VSS sg13g2_FILL8
XSTDFILL85_968 VDD VSS sg13g2_FILL8
XSTDFILL85_976 VDD VSS sg13g2_FILL8
XSTDFILL85_984 VDD VSS sg13g2_FILL8
XSTDFILL85_992 VDD VSS sg13g2_FILL8
XSTDFILL85_1000 VDD VSS sg13g2_FILL8
XSTDFILL85_1008 VDD VSS sg13g2_FILL8
XSTDFILL85_1016 VDD VSS sg13g2_FILL8
XSTDFILL85_1024 VDD VSS sg13g2_FILL8
XSTDFILL85_1032 VDD VSS sg13g2_FILL8
XSTDFILL85_1040 VDD VSS sg13g2_FILL8
XSTDFILL85_1048 VDD VSS sg13g2_FILL8
XSTDFILL85_1056 VDD VSS sg13g2_FILL8
XSTDFILL85_1064 VDD VSS sg13g2_FILL8
XSTDFILL85_1072 VDD VSS sg13g2_FILL8
XSTDFILL85_1080 VDD VSS sg13g2_FILL8
XSTDFILL85_1088 VDD VSS sg13g2_FILL8
XSTDFILL85_1096 VDD VSS sg13g2_FILL8
XSTDFILL85_1104 VDD VSS sg13g2_FILL8
XSTDFILL85_1112 VDD VSS sg13g2_FILL8
XSTDFILL85_1120 VDD VSS sg13g2_FILL8
XSTDFILL85_1128 VDD VSS sg13g2_FILL8
XSTDFILL85_1136 VDD VSS sg13g2_FILL8
XSTDFILL85_1144 VDD VSS sg13g2_FILL8
XSTDFILL85_1152 VDD VSS sg13g2_FILL8
XSTDFILL85_1160 VDD VSS sg13g2_FILL8
XSTDFILL85_1168 VDD VSS sg13g2_FILL8
XSTDFILL85_1176 VDD VSS sg13g2_FILL8
XSTDFILL85_1184 VDD VSS sg13g2_FILL8
XSTDFILL85_1192 VDD VSS sg13g2_FILL8
XSTDFILL85_1200 VDD VSS sg13g2_FILL8
XSTDFILL85_1208 VDD VSS sg13g2_FILL8
XSTDFILL85_1216 VDD VSS sg13g2_FILL8
XSTDFILL85_1224 VDD VSS sg13g2_FILL8
XSTDFILL85_1232 VDD VSS sg13g2_FILL8
XSTDFILL85_1240 VDD VSS sg13g2_FILL8
XSTDFILL85_1248 VDD VSS sg13g2_FILL8
XSTDFILL85_1256 VDD VSS sg13g2_FILL8
XSTDFILL85_1264 VDD VSS sg13g2_FILL8
XSTDFILL85_1272 VDD VSS sg13g2_FILL8
XSTDFILL85_1280 VDD VSS sg13g2_FILL8
XSTDFILL85_1288 VDD VSS sg13g2_FILL8
XSTDFILL85_1296 VDD VSS sg13g2_FILL8
XSTDFILL85_1304 VDD VSS sg13g2_FILL8
XSTDFILL85_1312 VDD VSS sg13g2_FILL8
XSTDFILL85_1320 VDD VSS sg13g2_FILL8
XSTDFILL85_1328 VDD VSS sg13g2_FILL8
XSTDFILL85_1336 VDD VSS sg13g2_FILL8
XSTDFILL85_1344 VDD VSS sg13g2_FILL8
XSTDFILL85_1352 VDD VSS sg13g2_FILL8
XSTDFILL85_1360 VDD VSS sg13g2_FILL8
XSTDFILL85_1368 VDD VSS sg13g2_FILL8
XSTDFILL85_1376 VDD VSS sg13g2_FILL8
XSTDFILL85_1384 VDD VSS sg13g2_FILL8
XSTDFILL85_1392 VDD VSS sg13g2_FILL8
XSTDFILL85_1400 VDD VSS sg13g2_FILL8
XSTDFILL85_1408 VDD VSS sg13g2_FILL8
XSTDFILL85_1416 VDD VSS sg13g2_FILL8
XSTDFILL85_1424 VDD VSS sg13g2_FILL8
XSTDFILL85_1432 VDD VSS sg13g2_FILL8
XSTDFILL85_1440 VDD VSS sg13g2_FILL8
XSTDFILL85_1448 VDD VSS sg13g2_FILL8
XSTDFILL85_1456 VDD VSS sg13g2_FILL8
XSTDFILL85_1464 VDD VSS sg13g2_FILL8
XSTDFILL85_1472 VDD VSS sg13g2_FILL8
XSTDFILL85_1480 VDD VSS sg13g2_FILL8
XSTDFILL85_1488 VDD VSS sg13g2_FILL8
XSTDFILL85_1496 VDD VSS sg13g2_FILL8
XSTDFILL85_1504 VDD VSS sg13g2_FILL8
XSTDFILL85_1512 VDD VSS sg13g2_FILL8
XSTDFILL85_1520 VDD VSS sg13g2_FILL8
XSTDFILL85_1528 VDD VSS sg13g2_FILL2
XSTDFILL85_1530 VDD VSS sg13g2_FILL1
XSTDFILL86_0 VDD VSS sg13g2_FILL8
XSTDFILL86_8 VDD VSS sg13g2_FILL8
XSTDFILL86_16 VDD VSS sg13g2_FILL8
XSTDFILL86_24 VDD VSS sg13g2_FILL8
XSTDFILL86_32 VDD VSS sg13g2_FILL8
XSTDFILL86_40 VDD VSS sg13g2_FILL8
XSTDFILL86_48 VDD VSS sg13g2_FILL8
XSTDFILL86_56 VDD VSS sg13g2_FILL8
XSTDFILL86_64 VDD VSS sg13g2_FILL8
XSTDFILL86_72 VDD VSS sg13g2_FILL8
XSTDFILL86_80 VDD VSS sg13g2_FILL8
XSTDFILL86_88 VDD VSS sg13g2_FILL8
XSTDFILL86_96 VDD VSS sg13g2_FILL8
XSTDFILL86_104 VDD VSS sg13g2_FILL8
XSTDFILL86_112 VDD VSS sg13g2_FILL8
XSTDFILL86_120 VDD VSS sg13g2_FILL8
XSTDFILL86_128 VDD VSS sg13g2_FILL8
XSTDFILL86_136 VDD VSS sg13g2_FILL8
XSTDFILL86_144 VDD VSS sg13g2_FILL8
XSTDFILL86_152 VDD VSS sg13g2_FILL8
XSTDFILL86_160 VDD VSS sg13g2_FILL8
XSTDFILL86_168 VDD VSS sg13g2_FILL8
XSTDFILL86_176 VDD VSS sg13g2_FILL8
XSTDFILL86_184 VDD VSS sg13g2_FILL8
XSTDFILL86_192 VDD VSS sg13g2_FILL8
XSTDFILL86_200 VDD VSS sg13g2_FILL8
XSTDFILL86_208 VDD VSS sg13g2_FILL8
XSTDFILL86_216 VDD VSS sg13g2_FILL8
XSTDFILL86_224 VDD VSS sg13g2_FILL8
XSTDFILL86_232 VDD VSS sg13g2_FILL8
XSTDFILL86_240 VDD VSS sg13g2_FILL8
XSTDFILL86_248 VDD VSS sg13g2_FILL8
XSTDFILL86_256 VDD VSS sg13g2_FILL8
XSTDFILL86_264 VDD VSS sg13g2_FILL8
XSTDFILL86_272 VDD VSS sg13g2_FILL8
XSTDFILL86_280 VDD VSS sg13g2_FILL8
XSTDFILL86_288 VDD VSS sg13g2_FILL8
XSTDFILL86_296 VDD VSS sg13g2_FILL8
XSTDFILL86_304 VDD VSS sg13g2_FILL8
XSTDFILL86_312 VDD VSS sg13g2_FILL8
XSTDFILL86_320 VDD VSS sg13g2_FILL8
XSTDFILL86_328 VDD VSS sg13g2_FILL8
XSTDFILL86_336 VDD VSS sg13g2_FILL8
XSTDFILL86_344 VDD VSS sg13g2_FILL8
XSTDFILL86_352 VDD VSS sg13g2_FILL8
XSTDFILL86_360 VDD VSS sg13g2_FILL8
XSTDFILL86_368 VDD VSS sg13g2_FILL8
XSTDFILL86_376 VDD VSS sg13g2_FILL8
XSTDFILL86_384 VDD VSS sg13g2_FILL8
XSTDFILL86_392 VDD VSS sg13g2_FILL8
XSTDFILL86_400 VDD VSS sg13g2_FILL8
XSTDFILL86_408 VDD VSS sg13g2_FILL8
XSTDFILL86_416 VDD VSS sg13g2_FILL8
XSTDFILL86_424 VDD VSS sg13g2_FILL8
XSTDFILL86_432 VDD VSS sg13g2_FILL8
XSTDFILL86_440 VDD VSS sg13g2_FILL8
XSTDFILL86_448 VDD VSS sg13g2_FILL8
XSTDFILL86_456 VDD VSS sg13g2_FILL8
XSTDFILL86_464 VDD VSS sg13g2_FILL8
XSTDFILL86_472 VDD VSS sg13g2_FILL8
XSTDFILL86_480 VDD VSS sg13g2_FILL8
XSTDFILL86_488 VDD VSS sg13g2_FILL8
XSTDFILL86_496 VDD VSS sg13g2_FILL8
XSTDFILL86_504 VDD VSS sg13g2_FILL8
XSTDFILL86_512 VDD VSS sg13g2_FILL8
XSTDFILL86_520 VDD VSS sg13g2_FILL8
XSTDFILL86_528 VDD VSS sg13g2_FILL8
XSTDFILL86_536 VDD VSS sg13g2_FILL8
XSTDFILL86_544 VDD VSS sg13g2_FILL8
XSTDFILL86_552 VDD VSS sg13g2_FILL8
XSTDFILL86_560 VDD VSS sg13g2_FILL8
XSTDFILL86_568 VDD VSS sg13g2_FILL8
XSTDFILL86_576 VDD VSS sg13g2_FILL8
XSTDFILL86_584 VDD VSS sg13g2_FILL8
XSTDFILL86_592 VDD VSS sg13g2_FILL8
XSTDFILL86_600 VDD VSS sg13g2_FILL8
XSTDFILL86_608 VDD VSS sg13g2_FILL8
XSTDFILL86_616 VDD VSS sg13g2_FILL8
XSTDFILL86_624 VDD VSS sg13g2_FILL8
XSTDFILL86_632 VDD VSS sg13g2_FILL8
XSTDFILL86_640 VDD VSS sg13g2_FILL8
XSTDFILL86_648 VDD VSS sg13g2_FILL8
XSTDFILL86_656 VDD VSS sg13g2_FILL8
XSTDFILL86_664 VDD VSS sg13g2_FILL8
XSTDFILL86_672 VDD VSS sg13g2_FILL8
XSTDFILL86_680 VDD VSS sg13g2_FILL8
XSTDFILL86_688 VDD VSS sg13g2_FILL8
XSTDFILL86_696 VDD VSS sg13g2_FILL8
XSTDFILL86_704 VDD VSS sg13g2_FILL8
XSTDFILL86_712 VDD VSS sg13g2_FILL8
XSTDFILL86_720 VDD VSS sg13g2_FILL8
XSTDFILL86_728 VDD VSS sg13g2_FILL8
XSTDFILL86_736 VDD VSS sg13g2_FILL8
XSTDFILL86_744 VDD VSS sg13g2_FILL8
XSTDFILL86_752 VDD VSS sg13g2_FILL8
XSTDFILL86_760 VDD VSS sg13g2_FILL8
XSTDFILL86_768 VDD VSS sg13g2_FILL8
XSTDFILL86_776 VDD VSS sg13g2_FILL8
XSTDFILL86_784 VDD VSS sg13g2_FILL8
XSTDFILL86_792 VDD VSS sg13g2_FILL8
XSTDFILL86_800 VDD VSS sg13g2_FILL8
XSTDFILL86_808 VDD VSS sg13g2_FILL8
XSTDFILL86_816 VDD VSS sg13g2_FILL8
XSTDFILL86_824 VDD VSS sg13g2_FILL8
XSTDFILL86_832 VDD VSS sg13g2_FILL8
XSTDFILL86_840 VDD VSS sg13g2_FILL8
XSTDFILL86_848 VDD VSS sg13g2_FILL8
XSTDFILL86_856 VDD VSS sg13g2_FILL8
XSTDFILL86_864 VDD VSS sg13g2_FILL8
XSTDFILL86_872 VDD VSS sg13g2_FILL8
XSTDFILL86_880 VDD VSS sg13g2_FILL8
XSTDFILL86_888 VDD VSS sg13g2_FILL8
XSTDFILL86_896 VDD VSS sg13g2_FILL8
XSTDFILL86_904 VDD VSS sg13g2_FILL8
XSTDFILL86_912 VDD VSS sg13g2_FILL8
XSTDFILL86_920 VDD VSS sg13g2_FILL8
XSTDFILL86_928 VDD VSS sg13g2_FILL8
XSTDFILL86_936 VDD VSS sg13g2_FILL8
XSTDFILL86_944 VDD VSS sg13g2_FILL8
XSTDFILL86_952 VDD VSS sg13g2_FILL8
XSTDFILL86_960 VDD VSS sg13g2_FILL8
XSTDFILL86_968 VDD VSS sg13g2_FILL8
XSTDFILL86_976 VDD VSS sg13g2_FILL8
XSTDFILL86_984 VDD VSS sg13g2_FILL8
XSTDFILL86_992 VDD VSS sg13g2_FILL8
XSTDFILL86_1000 VDD VSS sg13g2_FILL8
XSTDFILL86_1008 VDD VSS sg13g2_FILL8
XSTDFILL86_1016 VDD VSS sg13g2_FILL8
XSTDFILL86_1024 VDD VSS sg13g2_FILL8
XSTDFILL86_1032 VDD VSS sg13g2_FILL8
XSTDFILL86_1040 VDD VSS sg13g2_FILL8
XSTDFILL86_1048 VDD VSS sg13g2_FILL8
XSTDFILL86_1056 VDD VSS sg13g2_FILL8
XSTDFILL86_1064 VDD VSS sg13g2_FILL8
XSTDFILL86_1072 VDD VSS sg13g2_FILL8
XSTDFILL86_1080 VDD VSS sg13g2_FILL8
XSTDFILL86_1088 VDD VSS sg13g2_FILL8
XSTDFILL86_1096 VDD VSS sg13g2_FILL8
XSTDFILL86_1104 VDD VSS sg13g2_FILL8
XSTDFILL86_1112 VDD VSS sg13g2_FILL8
XSTDFILL86_1120 VDD VSS sg13g2_FILL8
XSTDFILL86_1128 VDD VSS sg13g2_FILL8
XSTDFILL86_1136 VDD VSS sg13g2_FILL8
XSTDFILL86_1144 VDD VSS sg13g2_FILL8
XSTDFILL86_1152 VDD VSS sg13g2_FILL8
XSTDFILL86_1160 VDD VSS sg13g2_FILL8
XSTDFILL86_1168 VDD VSS sg13g2_FILL8
XSTDFILL86_1176 VDD VSS sg13g2_FILL8
XSTDFILL86_1184 VDD VSS sg13g2_FILL8
XSTDFILL86_1192 VDD VSS sg13g2_FILL8
XSTDFILL86_1200 VDD VSS sg13g2_FILL8
XSTDFILL86_1208 VDD VSS sg13g2_FILL8
XSTDFILL86_1216 VDD VSS sg13g2_FILL8
XSTDFILL86_1224 VDD VSS sg13g2_FILL8
XSTDFILL86_1232 VDD VSS sg13g2_FILL8
XSTDFILL86_1240 VDD VSS sg13g2_FILL8
XSTDFILL86_1248 VDD VSS sg13g2_FILL8
XSTDFILL86_1256 VDD VSS sg13g2_FILL8
XSTDFILL86_1264 VDD VSS sg13g2_FILL8
XSTDFILL86_1272 VDD VSS sg13g2_FILL8
XSTDFILL86_1280 VDD VSS sg13g2_FILL8
XSTDFILL86_1288 VDD VSS sg13g2_FILL8
XSTDFILL86_1296 VDD VSS sg13g2_FILL8
XSTDFILL86_1304 VDD VSS sg13g2_FILL8
XSTDFILL86_1312 VDD VSS sg13g2_FILL8
XSTDFILL86_1320 VDD VSS sg13g2_FILL8
XSTDFILL86_1328 VDD VSS sg13g2_FILL8
XSTDFILL86_1336 VDD VSS sg13g2_FILL8
XSTDFILL86_1344 VDD VSS sg13g2_FILL8
XSTDFILL86_1352 VDD VSS sg13g2_FILL8
XSTDFILL86_1360 VDD VSS sg13g2_FILL8
XSTDFILL86_1368 VDD VSS sg13g2_FILL8
XSTDFILL86_1376 VDD VSS sg13g2_FILL8
XSTDFILL86_1384 VDD VSS sg13g2_FILL8
XSTDFILL86_1392 VDD VSS sg13g2_FILL8
XSTDFILL86_1400 VDD VSS sg13g2_FILL8
XSTDFILL86_1408 VDD VSS sg13g2_FILL8
XSTDFILL86_1416 VDD VSS sg13g2_FILL8
XSTDFILL86_1424 VDD VSS sg13g2_FILL8
XSTDFILL86_1432 VDD VSS sg13g2_FILL8
XSTDFILL86_1440 VDD VSS sg13g2_FILL8
XSTDFILL86_1448 VDD VSS sg13g2_FILL8
XSTDFILL86_1456 VDD VSS sg13g2_FILL8
XSTDFILL86_1464 VDD VSS sg13g2_FILL8
XSTDFILL86_1472 VDD VSS sg13g2_FILL8
XSTDFILL86_1480 VDD VSS sg13g2_FILL8
XSTDFILL86_1488 VDD VSS sg13g2_FILL8
XSTDFILL86_1496 VDD VSS sg13g2_FILL8
XSTDFILL86_1504 VDD VSS sg13g2_FILL8
XSTDFILL86_1512 VDD VSS sg13g2_FILL8
XSTDFILL86_1520 VDD VSS sg13g2_FILL8
XSTDFILL86_1528 VDD VSS sg13g2_FILL2
XSTDFILL86_1530 VDD VSS sg13g2_FILL1
XSTDFILL87_0 VDD VSS sg13g2_FILL8
XSTDFILL87_8 VDD VSS sg13g2_FILL8
XSTDFILL87_16 VDD VSS sg13g2_FILL8
XSTDFILL87_24 VDD VSS sg13g2_FILL8
XSTDFILL87_32 VDD VSS sg13g2_FILL8
XSTDFILL87_40 VDD VSS sg13g2_FILL8
XSTDFILL87_48 VDD VSS sg13g2_FILL8
XSTDFILL87_56 VDD VSS sg13g2_FILL8
XSTDFILL87_64 VDD VSS sg13g2_FILL8
XSTDFILL87_72 VDD VSS sg13g2_FILL8
XSTDFILL87_80 VDD VSS sg13g2_FILL8
XSTDFILL87_88 VDD VSS sg13g2_FILL8
XSTDFILL87_96 VDD VSS sg13g2_FILL8
XSTDFILL87_104 VDD VSS sg13g2_FILL8
XSTDFILL87_112 VDD VSS sg13g2_FILL8
XSTDFILL87_120 VDD VSS sg13g2_FILL8
XSTDFILL87_128 VDD VSS sg13g2_FILL8
XSTDFILL87_136 VDD VSS sg13g2_FILL8
XSTDFILL87_144 VDD VSS sg13g2_FILL8
XSTDFILL87_152 VDD VSS sg13g2_FILL8
XSTDFILL87_160 VDD VSS sg13g2_FILL8
XSTDFILL87_168 VDD VSS sg13g2_FILL8
XSTDFILL87_176 VDD VSS sg13g2_FILL8
XSTDFILL87_184 VDD VSS sg13g2_FILL8
XSTDFILL87_192 VDD VSS sg13g2_FILL8
XSTDFILL87_200 VDD VSS sg13g2_FILL8
XSTDFILL87_208 VDD VSS sg13g2_FILL8
XSTDFILL87_216 VDD VSS sg13g2_FILL8
XSTDFILL87_224 VDD VSS sg13g2_FILL8
XSTDFILL87_232 VDD VSS sg13g2_FILL8
XSTDFILL87_240 VDD VSS sg13g2_FILL8
XSTDFILL87_248 VDD VSS sg13g2_FILL8
XSTDFILL87_256 VDD VSS sg13g2_FILL8
XSTDFILL87_264 VDD VSS sg13g2_FILL8
XSTDFILL87_272 VDD VSS sg13g2_FILL8
XSTDFILL87_280 VDD VSS sg13g2_FILL8
XSTDFILL87_288 VDD VSS sg13g2_FILL8
XSTDFILL87_296 VDD VSS sg13g2_FILL8
XSTDFILL87_304 VDD VSS sg13g2_FILL8
XSTDFILL87_312 VDD VSS sg13g2_FILL8
XSTDFILL87_320 VDD VSS sg13g2_FILL8
XSTDFILL87_328 VDD VSS sg13g2_FILL8
XSTDFILL87_336 VDD VSS sg13g2_FILL8
XSTDFILL87_344 VDD VSS sg13g2_FILL8
XSTDFILL87_352 VDD VSS sg13g2_FILL8
XSTDFILL87_360 VDD VSS sg13g2_FILL8
XSTDFILL87_368 VDD VSS sg13g2_FILL8
XSTDFILL87_376 VDD VSS sg13g2_FILL8
XSTDFILL87_384 VDD VSS sg13g2_FILL8
XSTDFILL87_392 VDD VSS sg13g2_FILL8
XSTDFILL87_400 VDD VSS sg13g2_FILL8
XSTDFILL87_408 VDD VSS sg13g2_FILL8
XSTDFILL87_416 VDD VSS sg13g2_FILL8
XSTDFILL87_424 VDD VSS sg13g2_FILL8
XSTDFILL87_432 VDD VSS sg13g2_FILL8
XSTDFILL87_440 VDD VSS sg13g2_FILL8
XSTDFILL87_448 VDD VSS sg13g2_FILL8
XSTDFILL87_456 VDD VSS sg13g2_FILL8
XSTDFILL87_464 VDD VSS sg13g2_FILL8
XSTDFILL87_472 VDD VSS sg13g2_FILL8
XSTDFILL87_480 VDD VSS sg13g2_FILL8
XSTDFILL87_488 VDD VSS sg13g2_FILL8
XSTDFILL87_496 VDD VSS sg13g2_FILL8
XSTDFILL87_504 VDD VSS sg13g2_FILL8
XSTDFILL87_512 VDD VSS sg13g2_FILL8
XSTDFILL87_520 VDD VSS sg13g2_FILL8
XSTDFILL87_528 VDD VSS sg13g2_FILL8
XSTDFILL87_536 VDD VSS sg13g2_FILL8
XSTDFILL87_544 VDD VSS sg13g2_FILL8
XSTDFILL87_552 VDD VSS sg13g2_FILL8
XSTDFILL87_560 VDD VSS sg13g2_FILL8
XSTDFILL87_568 VDD VSS sg13g2_FILL8
XSTDFILL87_576 VDD VSS sg13g2_FILL8
XSTDFILL87_584 VDD VSS sg13g2_FILL8
XSTDFILL87_592 VDD VSS sg13g2_FILL8
XSTDFILL87_600 VDD VSS sg13g2_FILL8
XSTDFILL87_608 VDD VSS sg13g2_FILL8
XSTDFILL87_616 VDD VSS sg13g2_FILL8
XSTDFILL87_624 VDD VSS sg13g2_FILL8
XSTDFILL87_632 VDD VSS sg13g2_FILL8
XSTDFILL87_640 VDD VSS sg13g2_FILL8
XSTDFILL87_648 VDD VSS sg13g2_FILL8
XSTDFILL87_656 VDD VSS sg13g2_FILL8
XSTDFILL87_664 VDD VSS sg13g2_FILL8
XSTDFILL87_672 VDD VSS sg13g2_FILL8
XSTDFILL87_680 VDD VSS sg13g2_FILL8
XSTDFILL87_688 VDD VSS sg13g2_FILL8
XSTDFILL87_696 VDD VSS sg13g2_FILL8
XSTDFILL87_704 VDD VSS sg13g2_FILL8
XSTDFILL87_712 VDD VSS sg13g2_FILL8
XSTDFILL87_720 VDD VSS sg13g2_FILL8
XSTDFILL87_728 VDD VSS sg13g2_FILL8
XSTDFILL87_736 VDD VSS sg13g2_FILL8
XSTDFILL87_744 VDD VSS sg13g2_FILL8
XSTDFILL87_752 VDD VSS sg13g2_FILL8
XSTDFILL87_760 VDD VSS sg13g2_FILL8
XSTDFILL87_768 VDD VSS sg13g2_FILL8
XSTDFILL87_776 VDD VSS sg13g2_FILL8
XSTDFILL87_784 VDD VSS sg13g2_FILL8
XSTDFILL87_792 VDD VSS sg13g2_FILL8
XSTDFILL87_800 VDD VSS sg13g2_FILL8
XSTDFILL87_808 VDD VSS sg13g2_FILL8
XSTDFILL87_816 VDD VSS sg13g2_FILL8
XSTDFILL87_824 VDD VSS sg13g2_FILL8
XSTDFILL87_832 VDD VSS sg13g2_FILL8
XSTDFILL87_840 VDD VSS sg13g2_FILL8
XSTDFILL87_848 VDD VSS sg13g2_FILL8
XSTDFILL87_856 VDD VSS sg13g2_FILL8
XSTDFILL87_864 VDD VSS sg13g2_FILL8
XSTDFILL87_872 VDD VSS sg13g2_FILL8
XSTDFILL87_880 VDD VSS sg13g2_FILL8
XSTDFILL87_888 VDD VSS sg13g2_FILL8
XSTDFILL87_896 VDD VSS sg13g2_FILL8
XSTDFILL87_904 VDD VSS sg13g2_FILL8
XSTDFILL87_912 VDD VSS sg13g2_FILL8
XSTDFILL87_920 VDD VSS sg13g2_FILL8
XSTDFILL87_928 VDD VSS sg13g2_FILL8
XSTDFILL87_936 VDD VSS sg13g2_FILL8
XSTDFILL87_944 VDD VSS sg13g2_FILL8
XSTDFILL87_952 VDD VSS sg13g2_FILL8
XSTDFILL87_960 VDD VSS sg13g2_FILL8
XSTDFILL87_968 VDD VSS sg13g2_FILL8
XSTDFILL87_976 VDD VSS sg13g2_FILL8
XSTDFILL87_984 VDD VSS sg13g2_FILL8
XSTDFILL87_992 VDD VSS sg13g2_FILL8
XSTDFILL87_1000 VDD VSS sg13g2_FILL8
XSTDFILL87_1008 VDD VSS sg13g2_FILL8
XSTDFILL87_1016 VDD VSS sg13g2_FILL8
XSTDFILL87_1024 VDD VSS sg13g2_FILL8
XSTDFILL87_1032 VDD VSS sg13g2_FILL8
XSTDFILL87_1040 VDD VSS sg13g2_FILL8
XSTDFILL87_1048 VDD VSS sg13g2_FILL8
XSTDFILL87_1056 VDD VSS sg13g2_FILL8
XSTDFILL87_1064 VDD VSS sg13g2_FILL8
XSTDFILL87_1072 VDD VSS sg13g2_FILL8
XSTDFILL87_1080 VDD VSS sg13g2_FILL8
XSTDFILL87_1088 VDD VSS sg13g2_FILL8
XSTDFILL87_1096 VDD VSS sg13g2_FILL8
XSTDFILL87_1104 VDD VSS sg13g2_FILL8
XSTDFILL87_1112 VDD VSS sg13g2_FILL8
XSTDFILL87_1120 VDD VSS sg13g2_FILL8
XSTDFILL87_1128 VDD VSS sg13g2_FILL8
XSTDFILL87_1136 VDD VSS sg13g2_FILL8
XSTDFILL87_1144 VDD VSS sg13g2_FILL8
XSTDFILL87_1152 VDD VSS sg13g2_FILL8
XSTDFILL87_1160 VDD VSS sg13g2_FILL8
XSTDFILL87_1168 VDD VSS sg13g2_FILL8
XSTDFILL87_1176 VDD VSS sg13g2_FILL8
XSTDFILL87_1184 VDD VSS sg13g2_FILL8
XSTDFILL87_1192 VDD VSS sg13g2_FILL8
XSTDFILL87_1200 VDD VSS sg13g2_FILL8
XSTDFILL87_1208 VDD VSS sg13g2_FILL8
XSTDFILL87_1216 VDD VSS sg13g2_FILL8
XSTDFILL87_1224 VDD VSS sg13g2_FILL8
XSTDFILL87_1232 VDD VSS sg13g2_FILL8
XSTDFILL87_1240 VDD VSS sg13g2_FILL8
XSTDFILL87_1248 VDD VSS sg13g2_FILL8
XSTDFILL87_1256 VDD VSS sg13g2_FILL8
XSTDFILL87_1264 VDD VSS sg13g2_FILL8
XSTDFILL87_1272 VDD VSS sg13g2_FILL8
XSTDFILL87_1280 VDD VSS sg13g2_FILL8
XSTDFILL87_1288 VDD VSS sg13g2_FILL8
XSTDFILL87_1296 VDD VSS sg13g2_FILL8
XSTDFILL87_1304 VDD VSS sg13g2_FILL8
XSTDFILL87_1312 VDD VSS sg13g2_FILL8
XSTDFILL87_1320 VDD VSS sg13g2_FILL8
XSTDFILL87_1328 VDD VSS sg13g2_FILL8
XSTDFILL87_1336 VDD VSS sg13g2_FILL8
XSTDFILL87_1344 VDD VSS sg13g2_FILL8
XSTDFILL87_1352 VDD VSS sg13g2_FILL8
XSTDFILL87_1360 VDD VSS sg13g2_FILL8
XSTDFILL87_1368 VDD VSS sg13g2_FILL8
XSTDFILL87_1376 VDD VSS sg13g2_FILL8
XSTDFILL87_1384 VDD VSS sg13g2_FILL8
XSTDFILL87_1392 VDD VSS sg13g2_FILL8
XSTDFILL87_1400 VDD VSS sg13g2_FILL8
XSTDFILL87_1408 VDD VSS sg13g2_FILL8
XSTDFILL87_1416 VDD VSS sg13g2_FILL8
XSTDFILL87_1424 VDD VSS sg13g2_FILL8
XSTDFILL87_1432 VDD VSS sg13g2_FILL8
XSTDFILL87_1440 VDD VSS sg13g2_FILL8
XSTDFILL87_1448 VDD VSS sg13g2_FILL8
XSTDFILL87_1456 VDD VSS sg13g2_FILL8
XSTDFILL87_1464 VDD VSS sg13g2_FILL8
XSTDFILL87_1472 VDD VSS sg13g2_FILL8
XSTDFILL87_1480 VDD VSS sg13g2_FILL8
XSTDFILL87_1488 VDD VSS sg13g2_FILL8
XSTDFILL87_1496 VDD VSS sg13g2_FILL8
XSTDFILL87_1504 VDD VSS sg13g2_FILL8
XSTDFILL87_1512 VDD VSS sg13g2_FILL8
XSTDFILL87_1520 VDD VSS sg13g2_FILL8
XSTDFILL87_1528 VDD VSS sg13g2_FILL2
XSTDFILL87_1530 VDD VSS sg13g2_FILL1
XSTDFILL88_0 VDD VSS sg13g2_FILL8
XSTDFILL88_8 VDD VSS sg13g2_FILL8
XSTDFILL88_16 VDD VSS sg13g2_FILL8
XSTDFILL88_24 VDD VSS sg13g2_FILL8
XSTDFILL88_32 VDD VSS sg13g2_FILL8
XSTDFILL88_40 VDD VSS sg13g2_FILL8
XSTDFILL88_48 VDD VSS sg13g2_FILL8
XSTDFILL88_56 VDD VSS sg13g2_FILL8
XSTDFILL88_64 VDD VSS sg13g2_FILL8
XSTDFILL88_72 VDD VSS sg13g2_FILL8
XSTDFILL88_80 VDD VSS sg13g2_FILL8
XSTDFILL88_88 VDD VSS sg13g2_FILL8
XSTDFILL88_96 VDD VSS sg13g2_FILL8
XSTDFILL88_104 VDD VSS sg13g2_FILL8
XSTDFILL88_112 VDD VSS sg13g2_FILL8
XSTDFILL88_120 VDD VSS sg13g2_FILL8
XSTDFILL88_128 VDD VSS sg13g2_FILL8
XSTDFILL88_136 VDD VSS sg13g2_FILL8
XSTDFILL88_144 VDD VSS sg13g2_FILL8
XSTDFILL88_152 VDD VSS sg13g2_FILL8
XSTDFILL88_160 VDD VSS sg13g2_FILL8
XSTDFILL88_168 VDD VSS sg13g2_FILL8
XSTDFILL88_176 VDD VSS sg13g2_FILL8
XSTDFILL88_184 VDD VSS sg13g2_FILL8
XSTDFILL88_192 VDD VSS sg13g2_FILL8
XSTDFILL88_200 VDD VSS sg13g2_FILL8
XSTDFILL88_208 VDD VSS sg13g2_FILL8
XSTDFILL88_216 VDD VSS sg13g2_FILL8
XSTDFILL88_224 VDD VSS sg13g2_FILL8
XSTDFILL88_232 VDD VSS sg13g2_FILL8
XSTDFILL88_240 VDD VSS sg13g2_FILL8
XSTDFILL88_248 VDD VSS sg13g2_FILL8
XSTDFILL88_256 VDD VSS sg13g2_FILL8
XSTDFILL88_264 VDD VSS sg13g2_FILL8
XSTDFILL88_272 VDD VSS sg13g2_FILL8
XSTDFILL88_280 VDD VSS sg13g2_FILL8
XSTDFILL88_288 VDD VSS sg13g2_FILL8
XSTDFILL88_296 VDD VSS sg13g2_FILL8
XSTDFILL88_304 VDD VSS sg13g2_FILL8
XSTDFILL88_312 VDD VSS sg13g2_FILL8
XSTDFILL88_320 VDD VSS sg13g2_FILL8
XSTDFILL88_328 VDD VSS sg13g2_FILL8
XSTDFILL88_336 VDD VSS sg13g2_FILL8
XSTDFILL88_344 VDD VSS sg13g2_FILL8
XSTDFILL88_352 VDD VSS sg13g2_FILL8
XSTDFILL88_360 VDD VSS sg13g2_FILL8
XSTDFILL88_368 VDD VSS sg13g2_FILL8
XSTDFILL88_376 VDD VSS sg13g2_FILL8
XSTDFILL88_384 VDD VSS sg13g2_FILL8
XSTDFILL88_392 VDD VSS sg13g2_FILL8
XSTDFILL88_400 VDD VSS sg13g2_FILL8
XSTDFILL88_408 VDD VSS sg13g2_FILL8
XSTDFILL88_416 VDD VSS sg13g2_FILL8
XSTDFILL88_424 VDD VSS sg13g2_FILL8
XSTDFILL88_432 VDD VSS sg13g2_FILL8
XSTDFILL88_440 VDD VSS sg13g2_FILL8
XSTDFILL88_448 VDD VSS sg13g2_FILL8
XSTDFILL88_456 VDD VSS sg13g2_FILL8
XSTDFILL88_464 VDD VSS sg13g2_FILL8
XSTDFILL88_472 VDD VSS sg13g2_FILL8
XSTDFILL88_480 VDD VSS sg13g2_FILL8
XSTDFILL88_488 VDD VSS sg13g2_FILL8
XSTDFILL88_496 VDD VSS sg13g2_FILL8
XSTDFILL88_504 VDD VSS sg13g2_FILL8
XSTDFILL88_512 VDD VSS sg13g2_FILL8
XSTDFILL88_520 VDD VSS sg13g2_FILL8
XSTDFILL88_528 VDD VSS sg13g2_FILL8
XSTDFILL88_536 VDD VSS sg13g2_FILL8
XSTDFILL88_544 VDD VSS sg13g2_FILL8
XSTDFILL88_552 VDD VSS sg13g2_FILL8
XSTDFILL88_560 VDD VSS sg13g2_FILL8
XSTDFILL88_568 VDD VSS sg13g2_FILL8
XSTDFILL88_576 VDD VSS sg13g2_FILL8
XSTDFILL88_584 VDD VSS sg13g2_FILL8
XSTDFILL88_592 VDD VSS sg13g2_FILL8
XSTDFILL88_600 VDD VSS sg13g2_FILL8
XSTDFILL88_608 VDD VSS sg13g2_FILL8
XSTDFILL88_616 VDD VSS sg13g2_FILL8
XSTDFILL88_624 VDD VSS sg13g2_FILL8
XSTDFILL88_632 VDD VSS sg13g2_FILL8
XSTDFILL88_640 VDD VSS sg13g2_FILL8
XSTDFILL88_648 VDD VSS sg13g2_FILL8
XSTDFILL88_656 VDD VSS sg13g2_FILL8
XSTDFILL88_664 VDD VSS sg13g2_FILL8
XSTDFILL88_672 VDD VSS sg13g2_FILL8
XSTDFILL88_680 VDD VSS sg13g2_FILL8
XSTDFILL88_688 VDD VSS sg13g2_FILL8
XSTDFILL88_696 VDD VSS sg13g2_FILL8
XSTDFILL88_704 VDD VSS sg13g2_FILL8
XSTDFILL88_712 VDD VSS sg13g2_FILL8
XSTDFILL88_720 VDD VSS sg13g2_FILL8
XSTDFILL88_728 VDD VSS sg13g2_FILL8
XSTDFILL88_736 VDD VSS sg13g2_FILL8
XSTDFILL88_744 VDD VSS sg13g2_FILL8
XSTDFILL88_752 VDD VSS sg13g2_FILL8
XSTDFILL88_760 VDD VSS sg13g2_FILL8
XSTDFILL88_768 VDD VSS sg13g2_FILL8
XSTDFILL88_776 VDD VSS sg13g2_FILL8
XSTDFILL88_784 VDD VSS sg13g2_FILL8
XSTDFILL88_792 VDD VSS sg13g2_FILL8
XSTDFILL88_800 VDD VSS sg13g2_FILL8
XSTDFILL88_808 VDD VSS sg13g2_FILL8
XSTDFILL88_816 VDD VSS sg13g2_FILL8
XSTDFILL88_824 VDD VSS sg13g2_FILL8
XSTDFILL88_832 VDD VSS sg13g2_FILL8
XSTDFILL88_840 VDD VSS sg13g2_FILL8
XSTDFILL88_848 VDD VSS sg13g2_FILL8
XSTDFILL88_856 VDD VSS sg13g2_FILL8
XSTDFILL88_864 VDD VSS sg13g2_FILL8
XSTDFILL88_872 VDD VSS sg13g2_FILL8
XSTDFILL88_880 VDD VSS sg13g2_FILL8
XSTDFILL88_888 VDD VSS sg13g2_FILL8
XSTDFILL88_896 VDD VSS sg13g2_FILL8
XSTDFILL88_904 VDD VSS sg13g2_FILL8
XSTDFILL88_912 VDD VSS sg13g2_FILL8
XSTDFILL88_920 VDD VSS sg13g2_FILL8
XSTDFILL88_928 VDD VSS sg13g2_FILL8
XSTDFILL88_936 VDD VSS sg13g2_FILL8
XSTDFILL88_944 VDD VSS sg13g2_FILL8
XSTDFILL88_952 VDD VSS sg13g2_FILL8
XSTDFILL88_960 VDD VSS sg13g2_FILL8
XSTDFILL88_968 VDD VSS sg13g2_FILL8
XSTDFILL88_976 VDD VSS sg13g2_FILL8
XSTDFILL88_984 VDD VSS sg13g2_FILL8
XSTDFILL88_992 VDD VSS sg13g2_FILL8
XSTDFILL88_1000 VDD VSS sg13g2_FILL8
XSTDFILL88_1008 VDD VSS sg13g2_FILL8
XSTDFILL88_1016 VDD VSS sg13g2_FILL8
XSTDFILL88_1024 VDD VSS sg13g2_FILL8
XSTDFILL88_1032 VDD VSS sg13g2_FILL8
XSTDFILL88_1040 VDD VSS sg13g2_FILL8
XSTDFILL88_1048 VDD VSS sg13g2_FILL8
XSTDFILL88_1056 VDD VSS sg13g2_FILL8
XSTDFILL88_1064 VDD VSS sg13g2_FILL8
XSTDFILL88_1072 VDD VSS sg13g2_FILL8
XSTDFILL88_1080 VDD VSS sg13g2_FILL8
XSTDFILL88_1088 VDD VSS sg13g2_FILL8
XSTDFILL88_1096 VDD VSS sg13g2_FILL8
XSTDFILL88_1104 VDD VSS sg13g2_FILL8
XSTDFILL88_1112 VDD VSS sg13g2_FILL8
XSTDFILL88_1120 VDD VSS sg13g2_FILL8
XSTDFILL88_1128 VDD VSS sg13g2_FILL8
XSTDFILL88_1136 VDD VSS sg13g2_FILL8
XSTDFILL88_1144 VDD VSS sg13g2_FILL8
XSTDFILL88_1152 VDD VSS sg13g2_FILL8
XSTDFILL88_1160 VDD VSS sg13g2_FILL8
XSTDFILL88_1168 VDD VSS sg13g2_FILL8
XSTDFILL88_1176 VDD VSS sg13g2_FILL8
XSTDFILL88_1184 VDD VSS sg13g2_FILL8
XSTDFILL88_1192 VDD VSS sg13g2_FILL8
XSTDFILL88_1200 VDD VSS sg13g2_FILL8
XSTDFILL88_1208 VDD VSS sg13g2_FILL8
XSTDFILL88_1216 VDD VSS sg13g2_FILL8
XSTDFILL88_1224 VDD VSS sg13g2_FILL8
XSTDFILL88_1232 VDD VSS sg13g2_FILL8
XSTDFILL88_1240 VDD VSS sg13g2_FILL8
XSTDFILL88_1248 VDD VSS sg13g2_FILL8
XSTDFILL88_1256 VDD VSS sg13g2_FILL8
XSTDFILL88_1264 VDD VSS sg13g2_FILL8
XSTDFILL88_1272 VDD VSS sg13g2_FILL8
XSTDFILL88_1280 VDD VSS sg13g2_FILL8
XSTDFILL88_1288 VDD VSS sg13g2_FILL8
XSTDFILL88_1296 VDD VSS sg13g2_FILL8
XSTDFILL88_1304 VDD VSS sg13g2_FILL8
XSTDFILL88_1312 VDD VSS sg13g2_FILL8
XSTDFILL88_1320 VDD VSS sg13g2_FILL8
XSTDFILL88_1328 VDD VSS sg13g2_FILL8
XSTDFILL88_1336 VDD VSS sg13g2_FILL8
XSTDFILL88_1344 VDD VSS sg13g2_FILL8
XSTDFILL88_1352 VDD VSS sg13g2_FILL8
XSTDFILL88_1360 VDD VSS sg13g2_FILL8
XSTDFILL88_1368 VDD VSS sg13g2_FILL8
XSTDFILL88_1376 VDD VSS sg13g2_FILL8
XSTDFILL88_1384 VDD VSS sg13g2_FILL8
XSTDFILL88_1392 VDD VSS sg13g2_FILL8
XSTDFILL88_1400 VDD VSS sg13g2_FILL8
XSTDFILL88_1408 VDD VSS sg13g2_FILL8
XSTDFILL88_1416 VDD VSS sg13g2_FILL8
XSTDFILL88_1424 VDD VSS sg13g2_FILL8
XSTDFILL88_1432 VDD VSS sg13g2_FILL8
XSTDFILL88_1440 VDD VSS sg13g2_FILL8
XSTDFILL88_1448 VDD VSS sg13g2_FILL8
XSTDFILL88_1456 VDD VSS sg13g2_FILL8
XSTDFILL88_1464 VDD VSS sg13g2_FILL8
XSTDFILL88_1472 VDD VSS sg13g2_FILL8
XSTDFILL88_1480 VDD VSS sg13g2_FILL8
XSTDFILL88_1488 VDD VSS sg13g2_FILL8
XSTDFILL88_1496 VDD VSS sg13g2_FILL8
XSTDFILL88_1504 VDD VSS sg13g2_FILL8
XSTDFILL88_1512 VDD VSS sg13g2_FILL8
XSTDFILL88_1520 VDD VSS sg13g2_FILL8
XSTDFILL88_1528 VDD VSS sg13g2_FILL2
XSTDFILL88_1530 VDD VSS sg13g2_FILL1
XSTDFILL89_0 VDD VSS sg13g2_FILL8
XSTDFILL89_8 VDD VSS sg13g2_FILL8
XSTDFILL89_16 VDD VSS sg13g2_FILL8
XSTDFILL89_24 VDD VSS sg13g2_FILL8
XSTDFILL89_32 VDD VSS sg13g2_FILL8
XSTDFILL89_40 VDD VSS sg13g2_FILL8
XSTDFILL89_48 VDD VSS sg13g2_FILL8
XSTDFILL89_56 VDD VSS sg13g2_FILL8
XSTDFILL89_64 VDD VSS sg13g2_FILL8
XSTDFILL89_72 VDD VSS sg13g2_FILL8
XSTDFILL89_80 VDD VSS sg13g2_FILL8
XSTDFILL89_88 VDD VSS sg13g2_FILL8
XSTDFILL89_96 VDD VSS sg13g2_FILL8
XSTDFILL89_104 VDD VSS sg13g2_FILL8
XSTDFILL89_112 VDD VSS sg13g2_FILL8
XSTDFILL89_120 VDD VSS sg13g2_FILL8
XSTDFILL89_128 VDD VSS sg13g2_FILL8
XSTDFILL89_136 VDD VSS sg13g2_FILL8
XSTDFILL89_144 VDD VSS sg13g2_FILL8
XSTDFILL89_152 VDD VSS sg13g2_FILL8
XSTDFILL89_160 VDD VSS sg13g2_FILL8
XSTDFILL89_168 VDD VSS sg13g2_FILL8
XSTDFILL89_176 VDD VSS sg13g2_FILL8
XSTDFILL89_184 VDD VSS sg13g2_FILL8
XSTDFILL89_192 VDD VSS sg13g2_FILL8
XSTDFILL89_200 VDD VSS sg13g2_FILL8
XSTDFILL89_208 VDD VSS sg13g2_FILL8
XSTDFILL89_216 VDD VSS sg13g2_FILL8
XSTDFILL89_224 VDD VSS sg13g2_FILL8
XSTDFILL89_232 VDD VSS sg13g2_FILL8
XSTDFILL89_240 VDD VSS sg13g2_FILL8
XSTDFILL89_248 VDD VSS sg13g2_FILL8
XSTDFILL89_256 VDD VSS sg13g2_FILL8
XSTDFILL89_264 VDD VSS sg13g2_FILL8
XSTDFILL89_272 VDD VSS sg13g2_FILL8
XSTDFILL89_280 VDD VSS sg13g2_FILL8
XSTDFILL89_288 VDD VSS sg13g2_FILL8
XSTDFILL89_296 VDD VSS sg13g2_FILL8
XSTDFILL89_304 VDD VSS sg13g2_FILL8
XSTDFILL89_312 VDD VSS sg13g2_FILL8
XSTDFILL89_320 VDD VSS sg13g2_FILL8
XSTDFILL89_328 VDD VSS sg13g2_FILL8
XSTDFILL89_336 VDD VSS sg13g2_FILL8
XSTDFILL89_344 VDD VSS sg13g2_FILL8
XSTDFILL89_352 VDD VSS sg13g2_FILL8
XSTDFILL89_360 VDD VSS sg13g2_FILL8
XSTDFILL89_368 VDD VSS sg13g2_FILL8
XSTDFILL89_376 VDD VSS sg13g2_FILL8
XSTDFILL89_384 VDD VSS sg13g2_FILL8
XSTDFILL89_392 VDD VSS sg13g2_FILL8
XSTDFILL89_400 VDD VSS sg13g2_FILL8
XSTDFILL89_408 VDD VSS sg13g2_FILL8
XSTDFILL89_416 VDD VSS sg13g2_FILL8
XSTDFILL89_424 VDD VSS sg13g2_FILL8
XSTDFILL89_432 VDD VSS sg13g2_FILL8
XSTDFILL89_440 VDD VSS sg13g2_FILL8
XSTDFILL89_448 VDD VSS sg13g2_FILL8
XSTDFILL89_456 VDD VSS sg13g2_FILL8
XSTDFILL89_464 VDD VSS sg13g2_FILL8
XSTDFILL89_472 VDD VSS sg13g2_FILL8
XSTDFILL89_480 VDD VSS sg13g2_FILL8
XSTDFILL89_488 VDD VSS sg13g2_FILL8
XSTDFILL89_496 VDD VSS sg13g2_FILL8
XSTDFILL89_504 VDD VSS sg13g2_FILL8
XSTDFILL89_512 VDD VSS sg13g2_FILL8
XSTDFILL89_520 VDD VSS sg13g2_FILL8
XSTDFILL89_528 VDD VSS sg13g2_FILL8
XSTDFILL89_536 VDD VSS sg13g2_FILL8
XSTDFILL89_544 VDD VSS sg13g2_FILL8
XSTDFILL89_552 VDD VSS sg13g2_FILL8
XSTDFILL89_560 VDD VSS sg13g2_FILL8
XSTDFILL89_568 VDD VSS sg13g2_FILL8
XSTDFILL89_576 VDD VSS sg13g2_FILL8
XSTDFILL89_584 VDD VSS sg13g2_FILL8
XSTDFILL89_592 VDD VSS sg13g2_FILL8
XSTDFILL89_600 VDD VSS sg13g2_FILL8
XSTDFILL89_608 VDD VSS sg13g2_FILL8
XSTDFILL89_616 VDD VSS sg13g2_FILL8
XSTDFILL89_624 VDD VSS sg13g2_FILL8
XSTDFILL89_632 VDD VSS sg13g2_FILL8
XSTDFILL89_640 VDD VSS sg13g2_FILL8
XSTDFILL89_648 VDD VSS sg13g2_FILL8
XSTDFILL89_656 VDD VSS sg13g2_FILL8
XSTDFILL89_664 VDD VSS sg13g2_FILL8
XSTDFILL89_672 VDD VSS sg13g2_FILL8
XSTDFILL89_680 VDD VSS sg13g2_FILL8
XSTDFILL89_688 VDD VSS sg13g2_FILL8
XSTDFILL89_696 VDD VSS sg13g2_FILL8
XSTDFILL89_704 VDD VSS sg13g2_FILL8
XSTDFILL89_712 VDD VSS sg13g2_FILL8
XSTDFILL89_720 VDD VSS sg13g2_FILL8
XSTDFILL89_728 VDD VSS sg13g2_FILL8
XSTDFILL89_736 VDD VSS sg13g2_FILL8
XSTDFILL89_744 VDD VSS sg13g2_FILL8
XSTDFILL89_752 VDD VSS sg13g2_FILL8
XSTDFILL89_760 VDD VSS sg13g2_FILL8
XSTDFILL89_768 VDD VSS sg13g2_FILL8
XSTDFILL89_776 VDD VSS sg13g2_FILL8
XSTDFILL89_784 VDD VSS sg13g2_FILL8
XSTDFILL89_792 VDD VSS sg13g2_FILL8
XSTDFILL89_800 VDD VSS sg13g2_FILL8
XSTDFILL89_808 VDD VSS sg13g2_FILL8
XSTDFILL89_816 VDD VSS sg13g2_FILL8
XSTDFILL89_824 VDD VSS sg13g2_FILL8
XSTDFILL89_832 VDD VSS sg13g2_FILL8
XSTDFILL89_840 VDD VSS sg13g2_FILL8
XSTDFILL89_848 VDD VSS sg13g2_FILL8
XSTDFILL89_856 VDD VSS sg13g2_FILL8
XSTDFILL89_864 VDD VSS sg13g2_FILL8
XSTDFILL89_872 VDD VSS sg13g2_FILL8
XSTDFILL89_880 VDD VSS sg13g2_FILL8
XSTDFILL89_888 VDD VSS sg13g2_FILL8
XSTDFILL89_896 VDD VSS sg13g2_FILL8
XSTDFILL89_904 VDD VSS sg13g2_FILL8
XSTDFILL89_912 VDD VSS sg13g2_FILL8
XSTDFILL89_920 VDD VSS sg13g2_FILL8
XSTDFILL89_928 VDD VSS sg13g2_FILL8
XSTDFILL89_936 VDD VSS sg13g2_FILL8
XSTDFILL89_944 VDD VSS sg13g2_FILL8
XSTDFILL89_952 VDD VSS sg13g2_FILL8
XSTDFILL89_960 VDD VSS sg13g2_FILL8
XSTDFILL89_968 VDD VSS sg13g2_FILL8
XSTDFILL89_976 VDD VSS sg13g2_FILL8
XSTDFILL89_984 VDD VSS sg13g2_FILL8
XSTDFILL89_992 VDD VSS sg13g2_FILL8
XSTDFILL89_1000 VDD VSS sg13g2_FILL8
XSTDFILL89_1008 VDD VSS sg13g2_FILL8
XSTDFILL89_1016 VDD VSS sg13g2_FILL8
XSTDFILL89_1024 VDD VSS sg13g2_FILL8
XSTDFILL89_1032 VDD VSS sg13g2_FILL8
XSTDFILL89_1040 VDD VSS sg13g2_FILL8
XSTDFILL89_1048 VDD VSS sg13g2_FILL8
XSTDFILL89_1056 VDD VSS sg13g2_FILL8
XSTDFILL89_1064 VDD VSS sg13g2_FILL8
XSTDFILL89_1072 VDD VSS sg13g2_FILL8
XSTDFILL89_1080 VDD VSS sg13g2_FILL8
XSTDFILL89_1088 VDD VSS sg13g2_FILL8
XSTDFILL89_1096 VDD VSS sg13g2_FILL8
XSTDFILL89_1104 VDD VSS sg13g2_FILL8
XSTDFILL89_1112 VDD VSS sg13g2_FILL8
XSTDFILL89_1120 VDD VSS sg13g2_FILL8
XSTDFILL89_1128 VDD VSS sg13g2_FILL8
XSTDFILL89_1136 VDD VSS sg13g2_FILL8
XSTDFILL89_1144 VDD VSS sg13g2_FILL8
XSTDFILL89_1152 VDD VSS sg13g2_FILL8
XSTDFILL89_1160 VDD VSS sg13g2_FILL8
XSTDFILL89_1168 VDD VSS sg13g2_FILL8
XSTDFILL89_1176 VDD VSS sg13g2_FILL8
XSTDFILL89_1184 VDD VSS sg13g2_FILL8
XSTDFILL89_1192 VDD VSS sg13g2_FILL8
XSTDFILL89_1200 VDD VSS sg13g2_FILL8
XSTDFILL89_1208 VDD VSS sg13g2_FILL8
XSTDFILL89_1216 VDD VSS sg13g2_FILL8
XSTDFILL89_1224 VDD VSS sg13g2_FILL8
XSTDFILL89_1232 VDD VSS sg13g2_FILL8
XSTDFILL89_1240 VDD VSS sg13g2_FILL8
XSTDFILL89_1248 VDD VSS sg13g2_FILL8
XSTDFILL89_1256 VDD VSS sg13g2_FILL8
XSTDFILL89_1264 VDD VSS sg13g2_FILL8
XSTDFILL89_1272 VDD VSS sg13g2_FILL8
XSTDFILL89_1280 VDD VSS sg13g2_FILL8
XSTDFILL89_1288 VDD VSS sg13g2_FILL8
XSTDFILL89_1296 VDD VSS sg13g2_FILL8
XSTDFILL89_1304 VDD VSS sg13g2_FILL8
XSTDFILL89_1312 VDD VSS sg13g2_FILL8
XSTDFILL89_1320 VDD VSS sg13g2_FILL8
XSTDFILL89_1328 VDD VSS sg13g2_FILL8
XSTDFILL89_1336 VDD VSS sg13g2_FILL8
XSTDFILL89_1344 VDD VSS sg13g2_FILL8
XSTDFILL89_1352 VDD VSS sg13g2_FILL8
XSTDFILL89_1360 VDD VSS sg13g2_FILL8
XSTDFILL89_1368 VDD VSS sg13g2_FILL8
XSTDFILL89_1376 VDD VSS sg13g2_FILL8
XSTDFILL89_1384 VDD VSS sg13g2_FILL8
XSTDFILL89_1392 VDD VSS sg13g2_FILL8
XSTDFILL89_1400 VDD VSS sg13g2_FILL8
XSTDFILL89_1408 VDD VSS sg13g2_FILL8
XSTDFILL89_1416 VDD VSS sg13g2_FILL8
XSTDFILL89_1424 VDD VSS sg13g2_FILL8
XSTDFILL89_1432 VDD VSS sg13g2_FILL8
XSTDFILL89_1440 VDD VSS sg13g2_FILL8
XSTDFILL89_1448 VDD VSS sg13g2_FILL8
XSTDFILL89_1456 VDD VSS sg13g2_FILL8
XSTDFILL89_1464 VDD VSS sg13g2_FILL8
XSTDFILL89_1472 VDD VSS sg13g2_FILL8
XSTDFILL89_1480 VDD VSS sg13g2_FILL8
XSTDFILL89_1488 VDD VSS sg13g2_FILL8
XSTDFILL89_1496 VDD VSS sg13g2_FILL8
XSTDFILL89_1504 VDD VSS sg13g2_FILL8
XSTDFILL89_1512 VDD VSS sg13g2_FILL8
XSTDFILL89_1520 VDD VSS sg13g2_FILL8
XSTDFILL89_1528 VDD VSS sg13g2_FILL2
XSTDFILL89_1530 VDD VSS sg13g2_FILL1
XSTDFILL90_0 VDD VSS sg13g2_FILL8
XSTDFILL90_8 VDD VSS sg13g2_FILL8
XSTDFILL90_16 VDD VSS sg13g2_FILL8
XSTDFILL90_24 VDD VSS sg13g2_FILL8
XSTDFILL90_32 VDD VSS sg13g2_FILL8
XSTDFILL90_40 VDD VSS sg13g2_FILL8
XSTDFILL90_48 VDD VSS sg13g2_FILL8
XSTDFILL90_56 VDD VSS sg13g2_FILL8
XSTDFILL90_64 VDD VSS sg13g2_FILL8
XSTDFILL90_72 VDD VSS sg13g2_FILL8
XSTDFILL90_80 VDD VSS sg13g2_FILL8
XSTDFILL90_88 VDD VSS sg13g2_FILL8
XSTDFILL90_96 VDD VSS sg13g2_FILL8
XSTDFILL90_104 VDD VSS sg13g2_FILL8
XSTDFILL90_112 VDD VSS sg13g2_FILL8
XSTDFILL90_120 VDD VSS sg13g2_FILL8
XSTDFILL90_128 VDD VSS sg13g2_FILL8
XSTDFILL90_136 VDD VSS sg13g2_FILL8
XSTDFILL90_144 VDD VSS sg13g2_FILL8
XSTDFILL90_152 VDD VSS sg13g2_FILL8
XSTDFILL90_160 VDD VSS sg13g2_FILL8
XSTDFILL90_168 VDD VSS sg13g2_FILL8
XSTDFILL90_176 VDD VSS sg13g2_FILL8
XSTDFILL90_184 VDD VSS sg13g2_FILL8
XSTDFILL90_192 VDD VSS sg13g2_FILL8
XSTDFILL90_200 VDD VSS sg13g2_FILL8
XSTDFILL90_208 VDD VSS sg13g2_FILL8
XSTDFILL90_216 VDD VSS sg13g2_FILL8
XSTDFILL90_224 VDD VSS sg13g2_FILL8
XSTDFILL90_232 VDD VSS sg13g2_FILL8
XSTDFILL90_240 VDD VSS sg13g2_FILL8
XSTDFILL90_248 VDD VSS sg13g2_FILL8
XSTDFILL90_256 VDD VSS sg13g2_FILL8
XSTDFILL90_264 VDD VSS sg13g2_FILL8
XSTDFILL90_272 VDD VSS sg13g2_FILL8
XSTDFILL90_280 VDD VSS sg13g2_FILL8
XSTDFILL90_288 VDD VSS sg13g2_FILL8
XSTDFILL90_296 VDD VSS sg13g2_FILL8
XSTDFILL90_304 VDD VSS sg13g2_FILL8
XSTDFILL90_312 VDD VSS sg13g2_FILL8
XSTDFILL90_320 VDD VSS sg13g2_FILL8
XSTDFILL90_328 VDD VSS sg13g2_FILL8
XSTDFILL90_336 VDD VSS sg13g2_FILL8
XSTDFILL90_344 VDD VSS sg13g2_FILL8
XSTDFILL90_352 VDD VSS sg13g2_FILL8
XSTDFILL90_360 VDD VSS sg13g2_FILL8
XSTDFILL90_368 VDD VSS sg13g2_FILL8
XSTDFILL90_376 VDD VSS sg13g2_FILL8
XSTDFILL90_384 VDD VSS sg13g2_FILL8
XSTDFILL90_392 VDD VSS sg13g2_FILL8
XSTDFILL90_400 VDD VSS sg13g2_FILL8
XSTDFILL90_408 VDD VSS sg13g2_FILL8
XSTDFILL90_416 VDD VSS sg13g2_FILL8
XSTDFILL90_424 VDD VSS sg13g2_FILL8
XSTDFILL90_432 VDD VSS sg13g2_FILL8
XSTDFILL90_440 VDD VSS sg13g2_FILL8
XSTDFILL90_448 VDD VSS sg13g2_FILL8
XSTDFILL90_456 VDD VSS sg13g2_FILL8
XSTDFILL90_464 VDD VSS sg13g2_FILL8
XSTDFILL90_472 VDD VSS sg13g2_FILL8
XSTDFILL90_480 VDD VSS sg13g2_FILL8
XSTDFILL90_488 VDD VSS sg13g2_FILL8
XSTDFILL90_496 VDD VSS sg13g2_FILL8
XSTDFILL90_504 VDD VSS sg13g2_FILL8
XSTDFILL90_512 VDD VSS sg13g2_FILL8
XSTDFILL90_520 VDD VSS sg13g2_FILL8
XSTDFILL90_528 VDD VSS sg13g2_FILL8
XSTDFILL90_536 VDD VSS sg13g2_FILL8
XSTDFILL90_544 VDD VSS sg13g2_FILL8
XSTDFILL90_552 VDD VSS sg13g2_FILL8
XSTDFILL90_560 VDD VSS sg13g2_FILL8
XSTDFILL90_568 VDD VSS sg13g2_FILL8
XSTDFILL90_576 VDD VSS sg13g2_FILL8
XSTDFILL90_584 VDD VSS sg13g2_FILL8
XSTDFILL90_592 VDD VSS sg13g2_FILL8
XSTDFILL90_600 VDD VSS sg13g2_FILL8
XSTDFILL90_608 VDD VSS sg13g2_FILL8
XSTDFILL90_616 VDD VSS sg13g2_FILL8
XSTDFILL90_624 VDD VSS sg13g2_FILL8
XSTDFILL90_632 VDD VSS sg13g2_FILL8
XSTDFILL90_640 VDD VSS sg13g2_FILL8
XSTDFILL90_648 VDD VSS sg13g2_FILL8
XSTDFILL90_656 VDD VSS sg13g2_FILL8
XSTDFILL90_664 VDD VSS sg13g2_FILL8
XSTDFILL90_672 VDD VSS sg13g2_FILL8
XSTDFILL90_680 VDD VSS sg13g2_FILL8
XSTDFILL90_688 VDD VSS sg13g2_FILL8
XSTDFILL90_696 VDD VSS sg13g2_FILL8
XSTDFILL90_704 VDD VSS sg13g2_FILL8
XSTDFILL90_712 VDD VSS sg13g2_FILL8
XSTDFILL90_720 VDD VSS sg13g2_FILL8
XSTDFILL90_728 VDD VSS sg13g2_FILL8
XSTDFILL90_736 VDD VSS sg13g2_FILL8
XSTDFILL90_744 VDD VSS sg13g2_FILL8
XSTDFILL90_752 VDD VSS sg13g2_FILL8
XSTDFILL90_760 VDD VSS sg13g2_FILL8
XSTDFILL90_768 VDD VSS sg13g2_FILL8
XSTDFILL90_776 VDD VSS sg13g2_FILL8
XSTDFILL90_784 VDD VSS sg13g2_FILL8
XSTDFILL90_792 VDD VSS sg13g2_FILL8
XSTDFILL90_800 VDD VSS sg13g2_FILL8
XSTDFILL90_808 VDD VSS sg13g2_FILL8
XSTDFILL90_816 VDD VSS sg13g2_FILL8
XSTDFILL90_824 VDD VSS sg13g2_FILL8
XSTDFILL90_832 VDD VSS sg13g2_FILL8
XSTDFILL90_840 VDD VSS sg13g2_FILL8
XSTDFILL90_848 VDD VSS sg13g2_FILL8
XSTDFILL90_856 VDD VSS sg13g2_FILL8
XSTDFILL90_864 VDD VSS sg13g2_FILL8
XSTDFILL90_872 VDD VSS sg13g2_FILL8
XSTDFILL90_880 VDD VSS sg13g2_FILL8
XSTDFILL90_888 VDD VSS sg13g2_FILL8
XSTDFILL90_896 VDD VSS sg13g2_FILL8
XSTDFILL90_904 VDD VSS sg13g2_FILL8
XSTDFILL90_912 VDD VSS sg13g2_FILL8
XSTDFILL90_920 VDD VSS sg13g2_FILL8
XSTDFILL90_928 VDD VSS sg13g2_FILL8
XSTDFILL90_936 VDD VSS sg13g2_FILL8
XSTDFILL90_944 VDD VSS sg13g2_FILL8
XSTDFILL90_952 VDD VSS sg13g2_FILL8
XSTDFILL90_960 VDD VSS sg13g2_FILL8
XSTDFILL90_968 VDD VSS sg13g2_FILL8
XSTDFILL90_976 VDD VSS sg13g2_FILL8
XSTDFILL90_984 VDD VSS sg13g2_FILL8
XSTDFILL90_992 VDD VSS sg13g2_FILL8
XSTDFILL90_1000 VDD VSS sg13g2_FILL8
XSTDFILL90_1008 VDD VSS sg13g2_FILL8
XSTDFILL90_1016 VDD VSS sg13g2_FILL8
XSTDFILL90_1024 VDD VSS sg13g2_FILL8
XSTDFILL90_1032 VDD VSS sg13g2_FILL8
XSTDFILL90_1040 VDD VSS sg13g2_FILL8
XSTDFILL90_1048 VDD VSS sg13g2_FILL8
XSTDFILL90_1056 VDD VSS sg13g2_FILL8
XSTDFILL90_1064 VDD VSS sg13g2_FILL8
XSTDFILL90_1072 VDD VSS sg13g2_FILL8
XSTDFILL90_1080 VDD VSS sg13g2_FILL8
XSTDFILL90_1088 VDD VSS sg13g2_FILL8
XSTDFILL90_1096 VDD VSS sg13g2_FILL8
XSTDFILL90_1104 VDD VSS sg13g2_FILL8
XSTDFILL90_1112 VDD VSS sg13g2_FILL8
XSTDFILL90_1120 VDD VSS sg13g2_FILL8
XSTDFILL90_1128 VDD VSS sg13g2_FILL8
XSTDFILL90_1136 VDD VSS sg13g2_FILL8
XSTDFILL90_1144 VDD VSS sg13g2_FILL8
XSTDFILL90_1152 VDD VSS sg13g2_FILL8
XSTDFILL90_1160 VDD VSS sg13g2_FILL8
XSTDFILL90_1168 VDD VSS sg13g2_FILL8
XSTDFILL90_1176 VDD VSS sg13g2_FILL8
XSTDFILL90_1184 VDD VSS sg13g2_FILL8
XSTDFILL90_1192 VDD VSS sg13g2_FILL8
XSTDFILL90_1200 VDD VSS sg13g2_FILL8
XSTDFILL90_1208 VDD VSS sg13g2_FILL8
XSTDFILL90_1216 VDD VSS sg13g2_FILL8
XSTDFILL90_1224 VDD VSS sg13g2_FILL8
XSTDFILL90_1232 VDD VSS sg13g2_FILL8
XSTDFILL90_1240 VDD VSS sg13g2_FILL8
XSTDFILL90_1248 VDD VSS sg13g2_FILL8
XSTDFILL90_1256 VDD VSS sg13g2_FILL8
XSTDFILL90_1264 VDD VSS sg13g2_FILL8
XSTDFILL90_1272 VDD VSS sg13g2_FILL8
XSTDFILL90_1280 VDD VSS sg13g2_FILL8
XSTDFILL90_1288 VDD VSS sg13g2_FILL8
XSTDFILL90_1296 VDD VSS sg13g2_FILL8
XSTDFILL90_1304 VDD VSS sg13g2_FILL8
XSTDFILL90_1312 VDD VSS sg13g2_FILL8
XSTDFILL90_1320 VDD VSS sg13g2_FILL8
XSTDFILL90_1328 VDD VSS sg13g2_FILL8
XSTDFILL90_1336 VDD VSS sg13g2_FILL8
XSTDFILL90_1344 VDD VSS sg13g2_FILL8
XSTDFILL90_1352 VDD VSS sg13g2_FILL8
XSTDFILL90_1360 VDD VSS sg13g2_FILL8
XSTDFILL90_1368 VDD VSS sg13g2_FILL8
XSTDFILL90_1376 VDD VSS sg13g2_FILL8
XSTDFILL90_1384 VDD VSS sg13g2_FILL8
XSTDFILL90_1392 VDD VSS sg13g2_FILL8
XSTDFILL90_1400 VDD VSS sg13g2_FILL8
XSTDFILL90_1408 VDD VSS sg13g2_FILL8
XSTDFILL90_1416 VDD VSS sg13g2_FILL8
XSTDFILL90_1424 VDD VSS sg13g2_FILL8
XSTDFILL90_1432 VDD VSS sg13g2_FILL8
XSTDFILL90_1440 VDD VSS sg13g2_FILL8
XSTDFILL90_1448 VDD VSS sg13g2_FILL8
XSTDFILL90_1456 VDD VSS sg13g2_FILL8
XSTDFILL90_1464 VDD VSS sg13g2_FILL8
XSTDFILL90_1472 VDD VSS sg13g2_FILL8
XSTDFILL90_1480 VDD VSS sg13g2_FILL8
XSTDFILL90_1488 VDD VSS sg13g2_FILL8
XSTDFILL90_1496 VDD VSS sg13g2_FILL8
XSTDFILL90_1504 VDD VSS sg13g2_FILL8
XSTDFILL90_1512 VDD VSS sg13g2_FILL8
XSTDFILL90_1520 VDD VSS sg13g2_FILL8
XSTDFILL90_1528 VDD VSS sg13g2_FILL2
XSTDFILL90_1530 VDD VSS sg13g2_FILL1
XSTDFILL91_0 VDD VSS sg13g2_FILL8
XSTDFILL91_8 VDD VSS sg13g2_FILL8
XSTDFILL91_16 VDD VSS sg13g2_FILL8
XSTDFILL91_24 VDD VSS sg13g2_FILL8
XSTDFILL91_32 VDD VSS sg13g2_FILL8
XSTDFILL91_40 VDD VSS sg13g2_FILL8
XSTDFILL91_48 VDD VSS sg13g2_FILL8
XSTDFILL91_56 VDD VSS sg13g2_FILL8
XSTDFILL91_64 VDD VSS sg13g2_FILL8
XSTDFILL91_72 VDD VSS sg13g2_FILL8
XSTDFILL91_80 VDD VSS sg13g2_FILL8
XSTDFILL91_88 VDD VSS sg13g2_FILL8
XSTDFILL91_96 VDD VSS sg13g2_FILL8
XSTDFILL91_104 VDD VSS sg13g2_FILL8
XSTDFILL91_112 VDD VSS sg13g2_FILL8
XSTDFILL91_120 VDD VSS sg13g2_FILL8
XSTDFILL91_128 VDD VSS sg13g2_FILL8
XSTDFILL91_136 VDD VSS sg13g2_FILL8
XSTDFILL91_144 VDD VSS sg13g2_FILL8
XSTDFILL91_152 VDD VSS sg13g2_FILL8
XSTDFILL91_160 VDD VSS sg13g2_FILL8
XSTDFILL91_168 VDD VSS sg13g2_FILL8
XSTDFILL91_176 VDD VSS sg13g2_FILL8
XSTDFILL91_184 VDD VSS sg13g2_FILL8
XSTDFILL91_192 VDD VSS sg13g2_FILL8
XSTDFILL91_200 VDD VSS sg13g2_FILL8
XSTDFILL91_208 VDD VSS sg13g2_FILL8
XSTDFILL91_216 VDD VSS sg13g2_FILL8
XSTDFILL91_224 VDD VSS sg13g2_FILL8
XSTDFILL91_232 VDD VSS sg13g2_FILL8
XSTDFILL91_240 VDD VSS sg13g2_FILL8
XSTDFILL91_248 VDD VSS sg13g2_FILL8
XSTDFILL91_256 VDD VSS sg13g2_FILL8
XSTDFILL91_264 VDD VSS sg13g2_FILL8
XSTDFILL91_272 VDD VSS sg13g2_FILL8
XSTDFILL91_280 VDD VSS sg13g2_FILL8
XSTDFILL91_288 VDD VSS sg13g2_FILL8
XSTDFILL91_296 VDD VSS sg13g2_FILL8
XSTDFILL91_304 VDD VSS sg13g2_FILL8
XSTDFILL91_312 VDD VSS sg13g2_FILL8
XSTDFILL91_320 VDD VSS sg13g2_FILL8
XSTDFILL91_328 VDD VSS sg13g2_FILL8
XSTDFILL91_336 VDD VSS sg13g2_FILL8
XSTDFILL91_344 VDD VSS sg13g2_FILL8
XSTDFILL91_352 VDD VSS sg13g2_FILL8
XSTDFILL91_360 VDD VSS sg13g2_FILL8
XSTDFILL91_368 VDD VSS sg13g2_FILL8
XSTDFILL91_376 VDD VSS sg13g2_FILL8
XSTDFILL91_384 VDD VSS sg13g2_FILL8
XSTDFILL91_392 VDD VSS sg13g2_FILL8
XSTDFILL91_400 VDD VSS sg13g2_FILL8
XSTDFILL91_408 VDD VSS sg13g2_FILL8
XSTDFILL91_416 VDD VSS sg13g2_FILL8
XSTDFILL91_424 VDD VSS sg13g2_FILL8
XSTDFILL91_432 VDD VSS sg13g2_FILL8
XSTDFILL91_440 VDD VSS sg13g2_FILL8
XSTDFILL91_448 VDD VSS sg13g2_FILL8
XSTDFILL91_456 VDD VSS sg13g2_FILL8
XSTDFILL91_464 VDD VSS sg13g2_FILL8
XSTDFILL91_472 VDD VSS sg13g2_FILL8
XSTDFILL91_480 VDD VSS sg13g2_FILL8
XSTDFILL91_488 VDD VSS sg13g2_FILL8
XSTDFILL91_496 VDD VSS sg13g2_FILL8
XSTDFILL91_504 VDD VSS sg13g2_FILL8
XSTDFILL91_512 VDD VSS sg13g2_FILL8
XSTDFILL91_520 VDD VSS sg13g2_FILL8
XSTDFILL91_528 VDD VSS sg13g2_FILL8
XSTDFILL91_536 VDD VSS sg13g2_FILL8
XSTDFILL91_544 VDD VSS sg13g2_FILL8
XSTDFILL91_552 VDD VSS sg13g2_FILL8
XSTDFILL91_560 VDD VSS sg13g2_FILL8
XSTDFILL91_568 VDD VSS sg13g2_FILL8
XSTDFILL91_576 VDD VSS sg13g2_FILL8
XSTDFILL91_584 VDD VSS sg13g2_FILL8
XSTDFILL91_592 VDD VSS sg13g2_FILL8
XSTDFILL91_600 VDD VSS sg13g2_FILL8
XSTDFILL91_608 VDD VSS sg13g2_FILL8
XSTDFILL91_616 VDD VSS sg13g2_FILL8
XSTDFILL91_624 VDD VSS sg13g2_FILL8
XSTDFILL91_632 VDD VSS sg13g2_FILL8
XSTDFILL91_640 VDD VSS sg13g2_FILL8
XSTDFILL91_648 VDD VSS sg13g2_FILL8
XSTDFILL91_656 VDD VSS sg13g2_FILL8
XSTDFILL91_664 VDD VSS sg13g2_FILL8
XSTDFILL91_672 VDD VSS sg13g2_FILL8
XSTDFILL91_680 VDD VSS sg13g2_FILL8
XSTDFILL91_688 VDD VSS sg13g2_FILL8
XSTDFILL91_696 VDD VSS sg13g2_FILL8
XSTDFILL91_704 VDD VSS sg13g2_FILL8
XSTDFILL91_712 VDD VSS sg13g2_FILL8
XSTDFILL91_720 VDD VSS sg13g2_FILL8
XSTDFILL91_728 VDD VSS sg13g2_FILL8
XSTDFILL91_736 VDD VSS sg13g2_FILL8
XSTDFILL91_744 VDD VSS sg13g2_FILL8
XSTDFILL91_752 VDD VSS sg13g2_FILL8
XSTDFILL91_760 VDD VSS sg13g2_FILL8
XSTDFILL91_768 VDD VSS sg13g2_FILL8
XSTDFILL91_776 VDD VSS sg13g2_FILL8
XSTDFILL91_784 VDD VSS sg13g2_FILL8
XSTDFILL91_792 VDD VSS sg13g2_FILL8
XSTDFILL91_800 VDD VSS sg13g2_FILL8
XSTDFILL91_808 VDD VSS sg13g2_FILL8
XSTDFILL91_816 VDD VSS sg13g2_FILL8
XSTDFILL91_824 VDD VSS sg13g2_FILL8
XSTDFILL91_832 VDD VSS sg13g2_FILL8
XSTDFILL91_840 VDD VSS sg13g2_FILL8
XSTDFILL91_848 VDD VSS sg13g2_FILL8
XSTDFILL91_856 VDD VSS sg13g2_FILL8
XSTDFILL91_864 VDD VSS sg13g2_FILL8
XSTDFILL91_872 VDD VSS sg13g2_FILL8
XSTDFILL91_880 VDD VSS sg13g2_FILL8
XSTDFILL91_888 VDD VSS sg13g2_FILL8
XSTDFILL91_896 VDD VSS sg13g2_FILL8
XSTDFILL91_904 VDD VSS sg13g2_FILL8
XSTDFILL91_912 VDD VSS sg13g2_FILL8
XSTDFILL91_920 VDD VSS sg13g2_FILL8
XSTDFILL91_928 VDD VSS sg13g2_FILL8
XSTDFILL91_936 VDD VSS sg13g2_FILL8
XSTDFILL91_944 VDD VSS sg13g2_FILL8
XSTDFILL91_952 VDD VSS sg13g2_FILL8
XSTDFILL91_960 VDD VSS sg13g2_FILL8
XSTDFILL91_968 VDD VSS sg13g2_FILL8
XSTDFILL91_976 VDD VSS sg13g2_FILL8
XSTDFILL91_984 VDD VSS sg13g2_FILL8
XSTDFILL91_992 VDD VSS sg13g2_FILL8
XSTDFILL91_1000 VDD VSS sg13g2_FILL8
XSTDFILL91_1008 VDD VSS sg13g2_FILL8
XSTDFILL91_1016 VDD VSS sg13g2_FILL8
XSTDFILL91_1024 VDD VSS sg13g2_FILL8
XSTDFILL91_1032 VDD VSS sg13g2_FILL8
XSTDFILL91_1040 VDD VSS sg13g2_FILL8
XSTDFILL91_1048 VDD VSS sg13g2_FILL8
XSTDFILL91_1056 VDD VSS sg13g2_FILL8
XSTDFILL91_1064 VDD VSS sg13g2_FILL8
XSTDFILL91_1072 VDD VSS sg13g2_FILL8
XSTDFILL91_1080 VDD VSS sg13g2_FILL8
XSTDFILL91_1088 VDD VSS sg13g2_FILL8
XSTDFILL91_1096 VDD VSS sg13g2_FILL8
XSTDFILL91_1104 VDD VSS sg13g2_FILL8
XSTDFILL91_1112 VDD VSS sg13g2_FILL8
XSTDFILL91_1120 VDD VSS sg13g2_FILL8
XSTDFILL91_1128 VDD VSS sg13g2_FILL8
XSTDFILL91_1136 VDD VSS sg13g2_FILL8
XSTDFILL91_1144 VDD VSS sg13g2_FILL8
XSTDFILL91_1152 VDD VSS sg13g2_FILL8
XSTDFILL91_1160 VDD VSS sg13g2_FILL8
XSTDFILL91_1168 VDD VSS sg13g2_FILL8
XSTDFILL91_1176 VDD VSS sg13g2_FILL8
XSTDFILL91_1184 VDD VSS sg13g2_FILL8
XSTDFILL91_1192 VDD VSS sg13g2_FILL8
XSTDFILL91_1200 VDD VSS sg13g2_FILL8
XSTDFILL91_1208 VDD VSS sg13g2_FILL8
XSTDFILL91_1216 VDD VSS sg13g2_FILL8
XSTDFILL91_1224 VDD VSS sg13g2_FILL8
XSTDFILL91_1232 VDD VSS sg13g2_FILL8
XSTDFILL91_1240 VDD VSS sg13g2_FILL8
XSTDFILL91_1248 VDD VSS sg13g2_FILL8
XSTDFILL91_1256 VDD VSS sg13g2_FILL8
XSTDFILL91_1264 VDD VSS sg13g2_FILL8
XSTDFILL91_1272 VDD VSS sg13g2_FILL8
XSTDFILL91_1280 VDD VSS sg13g2_FILL8
XSTDFILL91_1288 VDD VSS sg13g2_FILL8
XSTDFILL91_1296 VDD VSS sg13g2_FILL8
XSTDFILL91_1304 VDD VSS sg13g2_FILL8
XSTDFILL91_1312 VDD VSS sg13g2_FILL8
XSTDFILL91_1320 VDD VSS sg13g2_FILL8
XSTDFILL91_1328 VDD VSS sg13g2_FILL8
XSTDFILL91_1336 VDD VSS sg13g2_FILL8
XSTDFILL91_1344 VDD VSS sg13g2_FILL8
XSTDFILL91_1352 VDD VSS sg13g2_FILL8
XSTDFILL91_1360 VDD VSS sg13g2_FILL8
XSTDFILL91_1368 VDD VSS sg13g2_FILL8
XSTDFILL91_1376 VDD VSS sg13g2_FILL8
XSTDFILL91_1384 VDD VSS sg13g2_FILL8
XSTDFILL91_1392 VDD VSS sg13g2_FILL8
XSTDFILL91_1400 VDD VSS sg13g2_FILL8
XSTDFILL91_1408 VDD VSS sg13g2_FILL8
XSTDFILL91_1416 VDD VSS sg13g2_FILL8
XSTDFILL91_1424 VDD VSS sg13g2_FILL8
XSTDFILL91_1432 VDD VSS sg13g2_FILL8
XSTDFILL91_1440 VDD VSS sg13g2_FILL8
XSTDFILL91_1448 VDD VSS sg13g2_FILL8
XSTDFILL91_1456 VDD VSS sg13g2_FILL8
XSTDFILL91_1464 VDD VSS sg13g2_FILL8
XSTDFILL91_1472 VDD VSS sg13g2_FILL8
XSTDFILL91_1480 VDD VSS sg13g2_FILL8
XSTDFILL91_1488 VDD VSS sg13g2_FILL8
XSTDFILL91_1496 VDD VSS sg13g2_FILL8
XSTDFILL91_1504 VDD VSS sg13g2_FILL8
XSTDFILL91_1512 VDD VSS sg13g2_FILL8
XSTDFILL91_1520 VDD VSS sg13g2_FILL8
XSTDFILL91_1528 VDD VSS sg13g2_FILL2
XSTDFILL91_1530 VDD VSS sg13g2_FILL1
XSTDFILL92_0 VDD VSS sg13g2_FILL8
XSTDFILL92_8 VDD VSS sg13g2_FILL8
XSTDFILL92_16 VDD VSS sg13g2_FILL8
XSTDFILL92_24 VDD VSS sg13g2_FILL8
XSTDFILL92_32 VDD VSS sg13g2_FILL8
XSTDFILL92_40 VDD VSS sg13g2_FILL8
XSTDFILL92_48 VDD VSS sg13g2_FILL8
XSTDFILL92_56 VDD VSS sg13g2_FILL8
XSTDFILL92_64 VDD VSS sg13g2_FILL8
XSTDFILL92_72 VDD VSS sg13g2_FILL8
XSTDFILL92_80 VDD VSS sg13g2_FILL8
XSTDFILL92_88 VDD VSS sg13g2_FILL8
XSTDFILL92_96 VDD VSS sg13g2_FILL8
XSTDFILL92_104 VDD VSS sg13g2_FILL8
XSTDFILL92_112 VDD VSS sg13g2_FILL8
XSTDFILL92_120 VDD VSS sg13g2_FILL8
XSTDFILL92_128 VDD VSS sg13g2_FILL8
XSTDFILL92_136 VDD VSS sg13g2_FILL8
XSTDFILL92_144 VDD VSS sg13g2_FILL8
XSTDFILL92_152 VDD VSS sg13g2_FILL8
XSTDFILL92_160 VDD VSS sg13g2_FILL8
XSTDFILL92_168 VDD VSS sg13g2_FILL8
XSTDFILL92_176 VDD VSS sg13g2_FILL8
XSTDFILL92_184 VDD VSS sg13g2_FILL8
XSTDFILL92_192 VDD VSS sg13g2_FILL8
XSTDFILL92_200 VDD VSS sg13g2_FILL8
XSTDFILL92_208 VDD VSS sg13g2_FILL8
XSTDFILL92_216 VDD VSS sg13g2_FILL8
XSTDFILL92_224 VDD VSS sg13g2_FILL8
XSTDFILL92_232 VDD VSS sg13g2_FILL8
XSTDFILL92_240 VDD VSS sg13g2_FILL8
XSTDFILL92_248 VDD VSS sg13g2_FILL8
XSTDFILL92_256 VDD VSS sg13g2_FILL8
XSTDFILL92_264 VDD VSS sg13g2_FILL8
XSTDFILL92_272 VDD VSS sg13g2_FILL8
XSTDFILL92_280 VDD VSS sg13g2_FILL8
XSTDFILL92_288 VDD VSS sg13g2_FILL8
XSTDFILL92_296 VDD VSS sg13g2_FILL8
XSTDFILL92_304 VDD VSS sg13g2_FILL8
XSTDFILL92_312 VDD VSS sg13g2_FILL8
XSTDFILL92_320 VDD VSS sg13g2_FILL8
XSTDFILL92_328 VDD VSS sg13g2_FILL8
XSTDFILL92_336 VDD VSS sg13g2_FILL8
XSTDFILL92_344 VDD VSS sg13g2_FILL8
XSTDFILL92_352 VDD VSS sg13g2_FILL8
XSTDFILL92_360 VDD VSS sg13g2_FILL8
XSTDFILL92_368 VDD VSS sg13g2_FILL8
XSTDFILL92_376 VDD VSS sg13g2_FILL8
XSTDFILL92_384 VDD VSS sg13g2_FILL8
XSTDFILL92_392 VDD VSS sg13g2_FILL8
XSTDFILL92_400 VDD VSS sg13g2_FILL8
XSTDFILL92_408 VDD VSS sg13g2_FILL8
XSTDFILL92_416 VDD VSS sg13g2_FILL8
XSTDFILL92_424 VDD VSS sg13g2_FILL8
XSTDFILL92_432 VDD VSS sg13g2_FILL8
XSTDFILL92_440 VDD VSS sg13g2_FILL8
XSTDFILL92_448 VDD VSS sg13g2_FILL8
XSTDFILL92_456 VDD VSS sg13g2_FILL8
XSTDFILL92_464 VDD VSS sg13g2_FILL8
XSTDFILL92_472 VDD VSS sg13g2_FILL8
XSTDFILL92_480 VDD VSS sg13g2_FILL8
XSTDFILL92_488 VDD VSS sg13g2_FILL8
XSTDFILL92_496 VDD VSS sg13g2_FILL8
XSTDFILL92_504 VDD VSS sg13g2_FILL8
XSTDFILL92_512 VDD VSS sg13g2_FILL8
XSTDFILL92_520 VDD VSS sg13g2_FILL8
XSTDFILL92_528 VDD VSS sg13g2_FILL8
XSTDFILL92_536 VDD VSS sg13g2_FILL8
XSTDFILL92_544 VDD VSS sg13g2_FILL8
XSTDFILL92_552 VDD VSS sg13g2_FILL8
XSTDFILL92_560 VDD VSS sg13g2_FILL8
XSTDFILL92_568 VDD VSS sg13g2_FILL8
XSTDFILL92_576 VDD VSS sg13g2_FILL8
XSTDFILL92_584 VDD VSS sg13g2_FILL8
XSTDFILL92_592 VDD VSS sg13g2_FILL8
XSTDFILL92_600 VDD VSS sg13g2_FILL8
XSTDFILL92_608 VDD VSS sg13g2_FILL8
XSTDFILL92_616 VDD VSS sg13g2_FILL8
XSTDFILL92_624 VDD VSS sg13g2_FILL8
XSTDFILL92_632 VDD VSS sg13g2_FILL8
XSTDFILL92_640 VDD VSS sg13g2_FILL8
XSTDFILL92_648 VDD VSS sg13g2_FILL8
XSTDFILL92_656 VDD VSS sg13g2_FILL8
XSTDFILL92_664 VDD VSS sg13g2_FILL8
XSTDFILL92_672 VDD VSS sg13g2_FILL8
XSTDFILL92_680 VDD VSS sg13g2_FILL8
XSTDFILL92_688 VDD VSS sg13g2_FILL8
XSTDFILL92_696 VDD VSS sg13g2_FILL8
XSTDFILL92_704 VDD VSS sg13g2_FILL8
XSTDFILL92_712 VDD VSS sg13g2_FILL8
XSTDFILL92_720 VDD VSS sg13g2_FILL8
XSTDFILL92_728 VDD VSS sg13g2_FILL8
XSTDFILL92_736 VDD VSS sg13g2_FILL8
XSTDFILL92_744 VDD VSS sg13g2_FILL8
XSTDFILL92_752 VDD VSS sg13g2_FILL8
XSTDFILL92_760 VDD VSS sg13g2_FILL8
XSTDFILL92_768 VDD VSS sg13g2_FILL8
XSTDFILL92_776 VDD VSS sg13g2_FILL8
XSTDFILL92_784 VDD VSS sg13g2_FILL8
XSTDFILL92_792 VDD VSS sg13g2_FILL8
XSTDFILL92_800 VDD VSS sg13g2_FILL8
XSTDFILL92_808 VDD VSS sg13g2_FILL8
XSTDFILL92_816 VDD VSS sg13g2_FILL8
XSTDFILL92_824 VDD VSS sg13g2_FILL8
XSTDFILL92_832 VDD VSS sg13g2_FILL8
XSTDFILL92_840 VDD VSS sg13g2_FILL8
XSTDFILL92_848 VDD VSS sg13g2_FILL8
XSTDFILL92_856 VDD VSS sg13g2_FILL8
XSTDFILL92_864 VDD VSS sg13g2_FILL8
XSTDFILL92_872 VDD VSS sg13g2_FILL8
XSTDFILL92_880 VDD VSS sg13g2_FILL8
XSTDFILL92_888 VDD VSS sg13g2_FILL8
XSTDFILL92_896 VDD VSS sg13g2_FILL8
XSTDFILL92_904 VDD VSS sg13g2_FILL8
XSTDFILL92_912 VDD VSS sg13g2_FILL8
XSTDFILL92_920 VDD VSS sg13g2_FILL8
XSTDFILL92_928 VDD VSS sg13g2_FILL8
XSTDFILL92_936 VDD VSS sg13g2_FILL8
XSTDFILL92_944 VDD VSS sg13g2_FILL8
XSTDFILL92_952 VDD VSS sg13g2_FILL8
XSTDFILL92_960 VDD VSS sg13g2_FILL8
XSTDFILL92_968 VDD VSS sg13g2_FILL8
XSTDFILL92_976 VDD VSS sg13g2_FILL8
XSTDFILL92_984 VDD VSS sg13g2_FILL8
XSTDFILL92_992 VDD VSS sg13g2_FILL8
XSTDFILL92_1000 VDD VSS sg13g2_FILL8
XSTDFILL92_1008 VDD VSS sg13g2_FILL8
XSTDFILL92_1016 VDD VSS sg13g2_FILL8
XSTDFILL92_1024 VDD VSS sg13g2_FILL8
XSTDFILL92_1032 VDD VSS sg13g2_FILL8
XSTDFILL92_1040 VDD VSS sg13g2_FILL8
XSTDFILL92_1048 VDD VSS sg13g2_FILL8
XSTDFILL92_1056 VDD VSS sg13g2_FILL8
XSTDFILL92_1064 VDD VSS sg13g2_FILL8
XSTDFILL92_1072 VDD VSS sg13g2_FILL8
XSTDFILL92_1080 VDD VSS sg13g2_FILL8
XSTDFILL92_1088 VDD VSS sg13g2_FILL8
XSTDFILL92_1096 VDD VSS sg13g2_FILL8
XSTDFILL92_1104 VDD VSS sg13g2_FILL8
XSTDFILL92_1112 VDD VSS sg13g2_FILL8
XSTDFILL92_1120 VDD VSS sg13g2_FILL8
XSTDFILL92_1128 VDD VSS sg13g2_FILL8
XSTDFILL92_1136 VDD VSS sg13g2_FILL8
XSTDFILL92_1144 VDD VSS sg13g2_FILL8
XSTDFILL92_1152 VDD VSS sg13g2_FILL8
XSTDFILL92_1160 VDD VSS sg13g2_FILL8
XSTDFILL92_1168 VDD VSS sg13g2_FILL8
XSTDFILL92_1176 VDD VSS sg13g2_FILL8
XSTDFILL92_1184 VDD VSS sg13g2_FILL8
XSTDFILL92_1192 VDD VSS sg13g2_FILL8
XSTDFILL92_1200 VDD VSS sg13g2_FILL8
XSTDFILL92_1208 VDD VSS sg13g2_FILL8
XSTDFILL92_1216 VDD VSS sg13g2_FILL8
XSTDFILL92_1224 VDD VSS sg13g2_FILL8
XSTDFILL92_1232 VDD VSS sg13g2_FILL8
XSTDFILL92_1240 VDD VSS sg13g2_FILL8
XSTDFILL92_1248 VDD VSS sg13g2_FILL8
XSTDFILL92_1256 VDD VSS sg13g2_FILL8
XSTDFILL92_1264 VDD VSS sg13g2_FILL8
XSTDFILL92_1272 VDD VSS sg13g2_FILL8
XSTDFILL92_1280 VDD VSS sg13g2_FILL8
XSTDFILL92_1288 VDD VSS sg13g2_FILL8
XSTDFILL92_1296 VDD VSS sg13g2_FILL8
XSTDFILL92_1304 VDD VSS sg13g2_FILL8
XSTDFILL92_1312 VDD VSS sg13g2_FILL8
XSTDFILL92_1320 VDD VSS sg13g2_FILL8
XSTDFILL92_1328 VDD VSS sg13g2_FILL8
XSTDFILL92_1336 VDD VSS sg13g2_FILL8
XSTDFILL92_1344 VDD VSS sg13g2_FILL8
XSTDFILL92_1352 VDD VSS sg13g2_FILL8
XSTDFILL92_1360 VDD VSS sg13g2_FILL8
XSTDFILL92_1368 VDD VSS sg13g2_FILL8
XSTDFILL92_1376 VDD VSS sg13g2_FILL8
XSTDFILL92_1384 VDD VSS sg13g2_FILL8
XSTDFILL92_1392 VDD VSS sg13g2_FILL8
XSTDFILL92_1400 VDD VSS sg13g2_FILL8
XSTDFILL92_1408 VDD VSS sg13g2_FILL8
XSTDFILL92_1416 VDD VSS sg13g2_FILL8
XSTDFILL92_1424 VDD VSS sg13g2_FILL8
XSTDFILL92_1432 VDD VSS sg13g2_FILL8
XSTDFILL92_1440 VDD VSS sg13g2_FILL8
XSTDFILL92_1448 VDD VSS sg13g2_FILL8
XSTDFILL92_1456 VDD VSS sg13g2_FILL8
XSTDFILL92_1464 VDD VSS sg13g2_FILL8
XSTDFILL92_1472 VDD VSS sg13g2_FILL8
XSTDFILL92_1480 VDD VSS sg13g2_FILL8
XSTDFILL92_1488 VDD VSS sg13g2_FILL8
XSTDFILL92_1496 VDD VSS sg13g2_FILL8
XSTDFILL92_1504 VDD VSS sg13g2_FILL8
XSTDFILL92_1512 VDD VSS sg13g2_FILL8
XSTDFILL92_1520 VDD VSS sg13g2_FILL8
XSTDFILL92_1528 VDD VSS sg13g2_FILL2
XSTDFILL92_1530 VDD VSS sg13g2_FILL1
XSTDFILL93_0 VDD VSS sg13g2_FILL8
XSTDFILL93_8 VDD VSS sg13g2_FILL8
XSTDFILL93_16 VDD VSS sg13g2_FILL8
XSTDFILL93_24 VDD VSS sg13g2_FILL8
XSTDFILL93_32 VDD VSS sg13g2_FILL8
XSTDFILL93_40 VDD VSS sg13g2_FILL8
XSTDFILL93_48 VDD VSS sg13g2_FILL8
XSTDFILL93_56 VDD VSS sg13g2_FILL8
XSTDFILL93_64 VDD VSS sg13g2_FILL8
XSTDFILL93_72 VDD VSS sg13g2_FILL8
XSTDFILL93_80 VDD VSS sg13g2_FILL8
XSTDFILL93_88 VDD VSS sg13g2_FILL8
XSTDFILL93_96 VDD VSS sg13g2_FILL8
XSTDFILL93_104 VDD VSS sg13g2_FILL8
XSTDFILL93_112 VDD VSS sg13g2_FILL8
XSTDFILL93_120 VDD VSS sg13g2_FILL8
XSTDFILL93_128 VDD VSS sg13g2_FILL8
XSTDFILL93_136 VDD VSS sg13g2_FILL8
XSTDFILL93_144 VDD VSS sg13g2_FILL8
XSTDFILL93_152 VDD VSS sg13g2_FILL8
XSTDFILL93_160 VDD VSS sg13g2_FILL8
XSTDFILL93_168 VDD VSS sg13g2_FILL8
XSTDFILL93_176 VDD VSS sg13g2_FILL8
XSTDFILL93_184 VDD VSS sg13g2_FILL8
XSTDFILL93_192 VDD VSS sg13g2_FILL8
XSTDFILL93_200 VDD VSS sg13g2_FILL8
XSTDFILL93_208 VDD VSS sg13g2_FILL8
XSTDFILL93_216 VDD VSS sg13g2_FILL8
XSTDFILL93_224 VDD VSS sg13g2_FILL8
XSTDFILL93_232 VDD VSS sg13g2_FILL8
XSTDFILL93_240 VDD VSS sg13g2_FILL8
XSTDFILL93_248 VDD VSS sg13g2_FILL8
XSTDFILL93_256 VDD VSS sg13g2_FILL8
XSTDFILL93_264 VDD VSS sg13g2_FILL8
XSTDFILL93_272 VDD VSS sg13g2_FILL8
XSTDFILL93_280 VDD VSS sg13g2_FILL8
XSTDFILL93_288 VDD VSS sg13g2_FILL8
XSTDFILL93_296 VDD VSS sg13g2_FILL8
XSTDFILL93_304 VDD VSS sg13g2_FILL8
XSTDFILL93_312 VDD VSS sg13g2_FILL8
XSTDFILL93_320 VDD VSS sg13g2_FILL8
XSTDFILL93_328 VDD VSS sg13g2_FILL8
XSTDFILL93_336 VDD VSS sg13g2_FILL8
XSTDFILL93_344 VDD VSS sg13g2_FILL8
XSTDFILL93_352 VDD VSS sg13g2_FILL8
XSTDFILL93_360 VDD VSS sg13g2_FILL8
XSTDFILL93_368 VDD VSS sg13g2_FILL8
XSTDFILL93_376 VDD VSS sg13g2_FILL8
XSTDFILL93_384 VDD VSS sg13g2_FILL8
XSTDFILL93_392 VDD VSS sg13g2_FILL8
XSTDFILL93_400 VDD VSS sg13g2_FILL8
XSTDFILL93_408 VDD VSS sg13g2_FILL8
XSTDFILL93_416 VDD VSS sg13g2_FILL8
XSTDFILL93_424 VDD VSS sg13g2_FILL8
XSTDFILL93_432 VDD VSS sg13g2_FILL8
XSTDFILL93_440 VDD VSS sg13g2_FILL8
XSTDFILL93_448 VDD VSS sg13g2_FILL8
XSTDFILL93_456 VDD VSS sg13g2_FILL8
XSTDFILL93_464 VDD VSS sg13g2_FILL8
XSTDFILL93_472 VDD VSS sg13g2_FILL8
XSTDFILL93_480 VDD VSS sg13g2_FILL8
XSTDFILL93_488 VDD VSS sg13g2_FILL8
XSTDFILL93_496 VDD VSS sg13g2_FILL8
XSTDFILL93_504 VDD VSS sg13g2_FILL8
XSTDFILL93_512 VDD VSS sg13g2_FILL8
XSTDFILL93_520 VDD VSS sg13g2_FILL8
XSTDFILL93_528 VDD VSS sg13g2_FILL8
XSTDFILL93_536 VDD VSS sg13g2_FILL8
XSTDFILL93_544 VDD VSS sg13g2_FILL8
XSTDFILL93_552 VDD VSS sg13g2_FILL8
XSTDFILL93_560 VDD VSS sg13g2_FILL8
XSTDFILL93_568 VDD VSS sg13g2_FILL8
XSTDFILL93_576 VDD VSS sg13g2_FILL8
XSTDFILL93_584 VDD VSS sg13g2_FILL8
XSTDFILL93_592 VDD VSS sg13g2_FILL8
XSTDFILL93_600 VDD VSS sg13g2_FILL8
XSTDFILL93_608 VDD VSS sg13g2_FILL8
XSTDFILL93_616 VDD VSS sg13g2_FILL8
XSTDFILL93_624 VDD VSS sg13g2_FILL8
XSTDFILL93_632 VDD VSS sg13g2_FILL8
XSTDFILL93_640 VDD VSS sg13g2_FILL8
XSTDFILL93_648 VDD VSS sg13g2_FILL8
XSTDFILL93_656 VDD VSS sg13g2_FILL8
XSTDFILL93_664 VDD VSS sg13g2_FILL8
XSTDFILL93_672 VDD VSS sg13g2_FILL8
XSTDFILL93_680 VDD VSS sg13g2_FILL8
XSTDFILL93_688 VDD VSS sg13g2_FILL8
XSTDFILL93_696 VDD VSS sg13g2_FILL8
XSTDFILL93_704 VDD VSS sg13g2_FILL8
XSTDFILL93_712 VDD VSS sg13g2_FILL8
XSTDFILL93_720 VDD VSS sg13g2_FILL8
XSTDFILL93_728 VDD VSS sg13g2_FILL8
XSTDFILL93_736 VDD VSS sg13g2_FILL8
XSTDFILL93_744 VDD VSS sg13g2_FILL8
XSTDFILL93_752 VDD VSS sg13g2_FILL8
XSTDFILL93_760 VDD VSS sg13g2_FILL8
XSTDFILL93_768 VDD VSS sg13g2_FILL8
XSTDFILL93_776 VDD VSS sg13g2_FILL8
XSTDFILL93_784 VDD VSS sg13g2_FILL8
XSTDFILL93_792 VDD VSS sg13g2_FILL8
XSTDFILL93_800 VDD VSS sg13g2_FILL8
XSTDFILL93_808 VDD VSS sg13g2_FILL8
XSTDFILL93_816 VDD VSS sg13g2_FILL8
XSTDFILL93_824 VDD VSS sg13g2_FILL8
XSTDFILL93_832 VDD VSS sg13g2_FILL8
XSTDFILL93_840 VDD VSS sg13g2_FILL8
XSTDFILL93_848 VDD VSS sg13g2_FILL8
XSTDFILL93_856 VDD VSS sg13g2_FILL8
XSTDFILL93_864 VDD VSS sg13g2_FILL8
XSTDFILL93_872 VDD VSS sg13g2_FILL8
XSTDFILL93_880 VDD VSS sg13g2_FILL8
XSTDFILL93_888 VDD VSS sg13g2_FILL8
XSTDFILL93_896 VDD VSS sg13g2_FILL8
XSTDFILL93_904 VDD VSS sg13g2_FILL8
XSTDFILL93_912 VDD VSS sg13g2_FILL8
XSTDFILL93_920 VDD VSS sg13g2_FILL8
XSTDFILL93_928 VDD VSS sg13g2_FILL8
XSTDFILL93_936 VDD VSS sg13g2_FILL8
XSTDFILL93_944 VDD VSS sg13g2_FILL8
XSTDFILL93_952 VDD VSS sg13g2_FILL8
XSTDFILL93_960 VDD VSS sg13g2_FILL8
XSTDFILL93_968 VDD VSS sg13g2_FILL8
XSTDFILL93_976 VDD VSS sg13g2_FILL8
XSTDFILL93_984 VDD VSS sg13g2_FILL8
XSTDFILL93_992 VDD VSS sg13g2_FILL8
XSTDFILL93_1000 VDD VSS sg13g2_FILL8
XSTDFILL93_1008 VDD VSS sg13g2_FILL8
XSTDFILL93_1016 VDD VSS sg13g2_FILL8
XSTDFILL93_1024 VDD VSS sg13g2_FILL8
XSTDFILL93_1032 VDD VSS sg13g2_FILL8
XSTDFILL93_1040 VDD VSS sg13g2_FILL8
XSTDFILL93_1048 VDD VSS sg13g2_FILL8
XSTDFILL93_1056 VDD VSS sg13g2_FILL8
XSTDFILL93_1064 VDD VSS sg13g2_FILL8
XSTDFILL93_1072 VDD VSS sg13g2_FILL8
XSTDFILL93_1080 VDD VSS sg13g2_FILL8
XSTDFILL93_1088 VDD VSS sg13g2_FILL8
XSTDFILL93_1096 VDD VSS sg13g2_FILL8
XSTDFILL93_1104 VDD VSS sg13g2_FILL8
XSTDFILL93_1112 VDD VSS sg13g2_FILL8
XSTDFILL93_1120 VDD VSS sg13g2_FILL8
XSTDFILL93_1128 VDD VSS sg13g2_FILL8
XSTDFILL93_1136 VDD VSS sg13g2_FILL8
XSTDFILL93_1144 VDD VSS sg13g2_FILL8
XSTDFILL93_1152 VDD VSS sg13g2_FILL8
XSTDFILL93_1160 VDD VSS sg13g2_FILL8
XSTDFILL93_1168 VDD VSS sg13g2_FILL8
XSTDFILL93_1176 VDD VSS sg13g2_FILL8
XSTDFILL93_1184 VDD VSS sg13g2_FILL8
XSTDFILL93_1192 VDD VSS sg13g2_FILL8
XSTDFILL93_1200 VDD VSS sg13g2_FILL8
XSTDFILL93_1208 VDD VSS sg13g2_FILL8
XSTDFILL93_1216 VDD VSS sg13g2_FILL8
XSTDFILL93_1224 VDD VSS sg13g2_FILL8
XSTDFILL93_1232 VDD VSS sg13g2_FILL8
XSTDFILL93_1240 VDD VSS sg13g2_FILL8
XSTDFILL93_1248 VDD VSS sg13g2_FILL8
XSTDFILL93_1256 VDD VSS sg13g2_FILL8
XSTDFILL93_1264 VDD VSS sg13g2_FILL8
XSTDFILL93_1272 VDD VSS sg13g2_FILL8
XSTDFILL93_1280 VDD VSS sg13g2_FILL8
XSTDFILL93_1288 VDD VSS sg13g2_FILL8
XSTDFILL93_1296 VDD VSS sg13g2_FILL8
XSTDFILL93_1304 VDD VSS sg13g2_FILL8
XSTDFILL93_1312 VDD VSS sg13g2_FILL8
XSTDFILL93_1320 VDD VSS sg13g2_FILL8
XSTDFILL93_1328 VDD VSS sg13g2_FILL8
XSTDFILL93_1336 VDD VSS sg13g2_FILL8
XSTDFILL93_1344 VDD VSS sg13g2_FILL8
XSTDFILL93_1352 VDD VSS sg13g2_FILL8
XSTDFILL93_1360 VDD VSS sg13g2_FILL8
XSTDFILL93_1368 VDD VSS sg13g2_FILL8
XSTDFILL93_1376 VDD VSS sg13g2_FILL8
XSTDFILL93_1384 VDD VSS sg13g2_FILL8
XSTDFILL93_1392 VDD VSS sg13g2_FILL8
XSTDFILL93_1400 VDD VSS sg13g2_FILL8
XSTDFILL93_1408 VDD VSS sg13g2_FILL8
XSTDFILL93_1416 VDD VSS sg13g2_FILL8
XSTDFILL93_1424 VDD VSS sg13g2_FILL8
XSTDFILL93_1432 VDD VSS sg13g2_FILL8
XSTDFILL93_1440 VDD VSS sg13g2_FILL8
XSTDFILL93_1448 VDD VSS sg13g2_FILL8
XSTDFILL93_1456 VDD VSS sg13g2_FILL8
XSTDFILL93_1464 VDD VSS sg13g2_FILL8
XSTDFILL93_1472 VDD VSS sg13g2_FILL8
XSTDFILL93_1480 VDD VSS sg13g2_FILL8
XSTDFILL93_1488 VDD VSS sg13g2_FILL8
XSTDFILL93_1496 VDD VSS sg13g2_FILL8
XSTDFILL93_1504 VDD VSS sg13g2_FILL8
XSTDFILL93_1512 VDD VSS sg13g2_FILL8
XSTDFILL93_1520 VDD VSS sg13g2_FILL8
XSTDFILL93_1528 VDD VSS sg13g2_FILL2
XSTDFILL93_1530 VDD VSS sg13g2_FILL1
XSTDFILL94_0 VDD VSS sg13g2_FILL8
XSTDFILL94_8 VDD VSS sg13g2_FILL8
XSTDFILL94_16 VDD VSS sg13g2_FILL8
XSTDFILL94_24 VDD VSS sg13g2_FILL8
XSTDFILL94_32 VDD VSS sg13g2_FILL8
XSTDFILL94_40 VDD VSS sg13g2_FILL8
XSTDFILL94_48 VDD VSS sg13g2_FILL8
XSTDFILL94_56 VDD VSS sg13g2_FILL8
XSTDFILL94_64 VDD VSS sg13g2_FILL8
XSTDFILL94_72 VDD VSS sg13g2_FILL8
XSTDFILL94_80 VDD VSS sg13g2_FILL8
XSTDFILL94_88 VDD VSS sg13g2_FILL8
XSTDFILL94_96 VDD VSS sg13g2_FILL8
XSTDFILL94_104 VDD VSS sg13g2_FILL8
XSTDFILL94_112 VDD VSS sg13g2_FILL8
XSTDFILL94_120 VDD VSS sg13g2_FILL8
XSTDFILL94_128 VDD VSS sg13g2_FILL8
XSTDFILL94_136 VDD VSS sg13g2_FILL8
XSTDFILL94_144 VDD VSS sg13g2_FILL8
XSTDFILL94_152 VDD VSS sg13g2_FILL8
XSTDFILL94_160 VDD VSS sg13g2_FILL8
XSTDFILL94_168 VDD VSS sg13g2_FILL8
XSTDFILL94_176 VDD VSS sg13g2_FILL8
XSTDFILL94_184 VDD VSS sg13g2_FILL8
XSTDFILL94_192 VDD VSS sg13g2_FILL8
XSTDFILL94_200 VDD VSS sg13g2_FILL8
XSTDFILL94_208 VDD VSS sg13g2_FILL8
XSTDFILL94_216 VDD VSS sg13g2_FILL8
XSTDFILL94_224 VDD VSS sg13g2_FILL8
XSTDFILL94_232 VDD VSS sg13g2_FILL8
XSTDFILL94_240 VDD VSS sg13g2_FILL8
XSTDFILL94_248 VDD VSS sg13g2_FILL8
XSTDFILL94_256 VDD VSS sg13g2_FILL8
XSTDFILL94_264 VDD VSS sg13g2_FILL8
XSTDFILL94_272 VDD VSS sg13g2_FILL8
XSTDFILL94_280 VDD VSS sg13g2_FILL8
XSTDFILL94_288 VDD VSS sg13g2_FILL8
XSTDFILL94_296 VDD VSS sg13g2_FILL8
XSTDFILL94_304 VDD VSS sg13g2_FILL8
XSTDFILL94_312 VDD VSS sg13g2_FILL8
XSTDFILL94_320 VDD VSS sg13g2_FILL8
XSTDFILL94_328 VDD VSS sg13g2_FILL8
XSTDFILL94_336 VDD VSS sg13g2_FILL8
XSTDFILL94_344 VDD VSS sg13g2_FILL8
XSTDFILL94_352 VDD VSS sg13g2_FILL8
XSTDFILL94_360 VDD VSS sg13g2_FILL8
XSTDFILL94_368 VDD VSS sg13g2_FILL8
XSTDFILL94_376 VDD VSS sg13g2_FILL8
XSTDFILL94_384 VDD VSS sg13g2_FILL8
XSTDFILL94_392 VDD VSS sg13g2_FILL8
XSTDFILL94_400 VDD VSS sg13g2_FILL8
XSTDFILL94_408 VDD VSS sg13g2_FILL8
XSTDFILL94_416 VDD VSS sg13g2_FILL8
XSTDFILL94_424 VDD VSS sg13g2_FILL8
XSTDFILL94_432 VDD VSS sg13g2_FILL8
XSTDFILL94_440 VDD VSS sg13g2_FILL8
XSTDFILL94_448 VDD VSS sg13g2_FILL8
XSTDFILL94_456 VDD VSS sg13g2_FILL8
XSTDFILL94_464 VDD VSS sg13g2_FILL8
XSTDFILL94_472 VDD VSS sg13g2_FILL8
XSTDFILL94_480 VDD VSS sg13g2_FILL8
XSTDFILL94_488 VDD VSS sg13g2_FILL8
XSTDFILL94_496 VDD VSS sg13g2_FILL8
XSTDFILL94_504 VDD VSS sg13g2_FILL8
XSTDFILL94_512 VDD VSS sg13g2_FILL8
XSTDFILL94_520 VDD VSS sg13g2_FILL8
XSTDFILL94_528 VDD VSS sg13g2_FILL8
XSTDFILL94_536 VDD VSS sg13g2_FILL8
XSTDFILL94_544 VDD VSS sg13g2_FILL8
XSTDFILL94_552 VDD VSS sg13g2_FILL8
XSTDFILL94_560 VDD VSS sg13g2_FILL8
XSTDFILL94_568 VDD VSS sg13g2_FILL8
XSTDFILL94_576 VDD VSS sg13g2_FILL8
XSTDFILL94_584 VDD VSS sg13g2_FILL8
XSTDFILL94_592 VDD VSS sg13g2_FILL8
XSTDFILL94_600 VDD VSS sg13g2_FILL8
XSTDFILL94_608 VDD VSS sg13g2_FILL8
XSTDFILL94_616 VDD VSS sg13g2_FILL8
XSTDFILL94_624 VDD VSS sg13g2_FILL8
XSTDFILL94_632 VDD VSS sg13g2_FILL8
XSTDFILL94_640 VDD VSS sg13g2_FILL8
XSTDFILL94_648 VDD VSS sg13g2_FILL8
XSTDFILL94_656 VDD VSS sg13g2_FILL8
XSTDFILL94_664 VDD VSS sg13g2_FILL8
XSTDFILL94_672 VDD VSS sg13g2_FILL8
XSTDFILL94_680 VDD VSS sg13g2_FILL8
XSTDFILL94_688 VDD VSS sg13g2_FILL8
XSTDFILL94_696 VDD VSS sg13g2_FILL8
XSTDFILL94_704 VDD VSS sg13g2_FILL8
XSTDFILL94_712 VDD VSS sg13g2_FILL8
XSTDFILL94_720 VDD VSS sg13g2_FILL8
XSTDFILL94_728 VDD VSS sg13g2_FILL8
XSTDFILL94_736 VDD VSS sg13g2_FILL8
XSTDFILL94_744 VDD VSS sg13g2_FILL8
XSTDFILL94_752 VDD VSS sg13g2_FILL8
XSTDFILL94_760 VDD VSS sg13g2_FILL8
XSTDFILL94_768 VDD VSS sg13g2_FILL8
XSTDFILL94_776 VDD VSS sg13g2_FILL8
XSTDFILL94_784 VDD VSS sg13g2_FILL8
XSTDFILL94_792 VDD VSS sg13g2_FILL8
XSTDFILL94_800 VDD VSS sg13g2_FILL8
XSTDFILL94_808 VDD VSS sg13g2_FILL8
XSTDFILL94_816 VDD VSS sg13g2_FILL8
XSTDFILL94_824 VDD VSS sg13g2_FILL8
XSTDFILL94_832 VDD VSS sg13g2_FILL8
XSTDFILL94_840 VDD VSS sg13g2_FILL8
XSTDFILL94_848 VDD VSS sg13g2_FILL8
XSTDFILL94_856 VDD VSS sg13g2_FILL8
XSTDFILL94_864 VDD VSS sg13g2_FILL8
XSTDFILL94_872 VDD VSS sg13g2_FILL8
XSTDFILL94_880 VDD VSS sg13g2_FILL8
XSTDFILL94_888 VDD VSS sg13g2_FILL8
XSTDFILL94_896 VDD VSS sg13g2_FILL8
XSTDFILL94_904 VDD VSS sg13g2_FILL8
XSTDFILL94_912 VDD VSS sg13g2_FILL8
XSTDFILL94_920 VDD VSS sg13g2_FILL8
XSTDFILL94_928 VDD VSS sg13g2_FILL8
XSTDFILL94_936 VDD VSS sg13g2_FILL8
XSTDFILL94_944 VDD VSS sg13g2_FILL8
XSTDFILL94_952 VDD VSS sg13g2_FILL8
XSTDFILL94_960 VDD VSS sg13g2_FILL8
XSTDFILL94_968 VDD VSS sg13g2_FILL8
XSTDFILL94_976 VDD VSS sg13g2_FILL8
XSTDFILL94_984 VDD VSS sg13g2_FILL8
XSTDFILL94_992 VDD VSS sg13g2_FILL8
XSTDFILL94_1000 VDD VSS sg13g2_FILL8
XSTDFILL94_1008 VDD VSS sg13g2_FILL8
XSTDFILL94_1016 VDD VSS sg13g2_FILL8
XSTDFILL94_1024 VDD VSS sg13g2_FILL8
XSTDFILL94_1032 VDD VSS sg13g2_FILL8
XSTDFILL94_1040 VDD VSS sg13g2_FILL8
XSTDFILL94_1048 VDD VSS sg13g2_FILL8
XSTDFILL94_1056 VDD VSS sg13g2_FILL8
XSTDFILL94_1064 VDD VSS sg13g2_FILL8
XSTDFILL94_1072 VDD VSS sg13g2_FILL8
XSTDFILL94_1080 VDD VSS sg13g2_FILL8
XSTDFILL94_1088 VDD VSS sg13g2_FILL8
XSTDFILL94_1096 VDD VSS sg13g2_FILL8
XSTDFILL94_1104 VDD VSS sg13g2_FILL8
XSTDFILL94_1112 VDD VSS sg13g2_FILL8
XSTDFILL94_1120 VDD VSS sg13g2_FILL8
XSTDFILL94_1128 VDD VSS sg13g2_FILL8
XSTDFILL94_1136 VDD VSS sg13g2_FILL8
XSTDFILL94_1144 VDD VSS sg13g2_FILL8
XSTDFILL94_1152 VDD VSS sg13g2_FILL8
XSTDFILL94_1160 VDD VSS sg13g2_FILL8
XSTDFILL94_1168 VDD VSS sg13g2_FILL8
XSTDFILL94_1176 VDD VSS sg13g2_FILL8
XSTDFILL94_1184 VDD VSS sg13g2_FILL8
XSTDFILL94_1192 VDD VSS sg13g2_FILL8
XSTDFILL94_1200 VDD VSS sg13g2_FILL8
XSTDFILL94_1208 VDD VSS sg13g2_FILL8
XSTDFILL94_1216 VDD VSS sg13g2_FILL8
XSTDFILL94_1224 VDD VSS sg13g2_FILL8
XSTDFILL94_1232 VDD VSS sg13g2_FILL8
XSTDFILL94_1240 VDD VSS sg13g2_FILL8
XSTDFILL94_1248 VDD VSS sg13g2_FILL8
XSTDFILL94_1256 VDD VSS sg13g2_FILL8
XSTDFILL94_1264 VDD VSS sg13g2_FILL8
XSTDFILL94_1272 VDD VSS sg13g2_FILL8
XSTDFILL94_1280 VDD VSS sg13g2_FILL8
XSTDFILL94_1288 VDD VSS sg13g2_FILL8
XSTDFILL94_1296 VDD VSS sg13g2_FILL8
XSTDFILL94_1304 VDD VSS sg13g2_FILL8
XSTDFILL94_1312 VDD VSS sg13g2_FILL8
XSTDFILL94_1320 VDD VSS sg13g2_FILL8
XSTDFILL94_1328 VDD VSS sg13g2_FILL8
XSTDFILL94_1336 VDD VSS sg13g2_FILL8
XSTDFILL94_1344 VDD VSS sg13g2_FILL8
XSTDFILL94_1352 VDD VSS sg13g2_FILL8
XSTDFILL94_1360 VDD VSS sg13g2_FILL8
XSTDFILL94_1368 VDD VSS sg13g2_FILL8
XSTDFILL94_1376 VDD VSS sg13g2_FILL8
XSTDFILL94_1384 VDD VSS sg13g2_FILL8
XSTDFILL94_1392 VDD VSS sg13g2_FILL8
XSTDFILL94_1400 VDD VSS sg13g2_FILL8
XSTDFILL94_1408 VDD VSS sg13g2_FILL8
XSTDFILL94_1416 VDD VSS sg13g2_FILL8
XSTDFILL94_1424 VDD VSS sg13g2_FILL8
XSTDFILL94_1432 VDD VSS sg13g2_FILL8
XSTDFILL94_1440 VDD VSS sg13g2_FILL8
XSTDFILL94_1448 VDD VSS sg13g2_FILL8
XSTDFILL94_1456 VDD VSS sg13g2_FILL8
XSTDFILL94_1464 VDD VSS sg13g2_FILL8
XSTDFILL94_1472 VDD VSS sg13g2_FILL8
XSTDFILL94_1480 VDD VSS sg13g2_FILL8
XSTDFILL94_1488 VDD VSS sg13g2_FILL8
XSTDFILL94_1496 VDD VSS sg13g2_FILL8
XSTDFILL94_1504 VDD VSS sg13g2_FILL8
XSTDFILL94_1512 VDD VSS sg13g2_FILL8
XSTDFILL94_1520 VDD VSS sg13g2_FILL8
XSTDFILL94_1528 VDD VSS sg13g2_FILL2
XSTDFILL94_1530 VDD VSS sg13g2_FILL1
XSTDFILL95_0 VDD VSS sg13g2_FILL8
XSTDFILL95_8 VDD VSS sg13g2_FILL8
XSTDFILL95_16 VDD VSS sg13g2_FILL8
XSTDFILL95_24 VDD VSS sg13g2_FILL8
XSTDFILL95_32 VDD VSS sg13g2_FILL8
XSTDFILL95_40 VDD VSS sg13g2_FILL8
XSTDFILL95_48 VDD VSS sg13g2_FILL8
XSTDFILL95_56 VDD VSS sg13g2_FILL8
XSTDFILL95_64 VDD VSS sg13g2_FILL8
XSTDFILL95_72 VDD VSS sg13g2_FILL8
XSTDFILL95_80 VDD VSS sg13g2_FILL8
XSTDFILL95_88 VDD VSS sg13g2_FILL8
XSTDFILL95_96 VDD VSS sg13g2_FILL8
XSTDFILL95_104 VDD VSS sg13g2_FILL8
XSTDFILL95_112 VDD VSS sg13g2_FILL8
XSTDFILL95_120 VDD VSS sg13g2_FILL8
XSTDFILL95_128 VDD VSS sg13g2_FILL8
XSTDFILL95_136 VDD VSS sg13g2_FILL8
XSTDFILL95_144 VDD VSS sg13g2_FILL8
XSTDFILL95_152 VDD VSS sg13g2_FILL8
XSTDFILL95_160 VDD VSS sg13g2_FILL8
XSTDFILL95_168 VDD VSS sg13g2_FILL8
XSTDFILL95_176 VDD VSS sg13g2_FILL8
XSTDFILL95_184 VDD VSS sg13g2_FILL8
XSTDFILL95_192 VDD VSS sg13g2_FILL8
XSTDFILL95_200 VDD VSS sg13g2_FILL8
XSTDFILL95_208 VDD VSS sg13g2_FILL8
XSTDFILL95_216 VDD VSS sg13g2_FILL8
XSTDFILL95_224 VDD VSS sg13g2_FILL8
XSTDFILL95_232 VDD VSS sg13g2_FILL8
XSTDFILL95_240 VDD VSS sg13g2_FILL8
XSTDFILL95_248 VDD VSS sg13g2_FILL8
XSTDFILL95_256 VDD VSS sg13g2_FILL8
XSTDFILL95_264 VDD VSS sg13g2_FILL8
XSTDFILL95_272 VDD VSS sg13g2_FILL8
XSTDFILL95_280 VDD VSS sg13g2_FILL8
XSTDFILL95_288 VDD VSS sg13g2_FILL8
XSTDFILL95_296 VDD VSS sg13g2_FILL8
XSTDFILL95_304 VDD VSS sg13g2_FILL8
XSTDFILL95_312 VDD VSS sg13g2_FILL8
XSTDFILL95_320 VDD VSS sg13g2_FILL8
XSTDFILL95_328 VDD VSS sg13g2_FILL8
XSTDFILL95_336 VDD VSS sg13g2_FILL8
XSTDFILL95_344 VDD VSS sg13g2_FILL8
XSTDFILL95_352 VDD VSS sg13g2_FILL8
XSTDFILL95_360 VDD VSS sg13g2_FILL8
XSTDFILL95_368 VDD VSS sg13g2_FILL8
XSTDFILL95_376 VDD VSS sg13g2_FILL8
XSTDFILL95_384 VDD VSS sg13g2_FILL8
XSTDFILL95_392 VDD VSS sg13g2_FILL8
XSTDFILL95_400 VDD VSS sg13g2_FILL8
XSTDFILL95_408 VDD VSS sg13g2_FILL8
XSTDFILL95_416 VDD VSS sg13g2_FILL8
XSTDFILL95_424 VDD VSS sg13g2_FILL8
XSTDFILL95_432 VDD VSS sg13g2_FILL8
XSTDFILL95_440 VDD VSS sg13g2_FILL8
XSTDFILL95_448 VDD VSS sg13g2_FILL8
XSTDFILL95_456 VDD VSS sg13g2_FILL8
XSTDFILL95_464 VDD VSS sg13g2_FILL8
XSTDFILL95_472 VDD VSS sg13g2_FILL8
XSTDFILL95_480 VDD VSS sg13g2_FILL8
XSTDFILL95_488 VDD VSS sg13g2_FILL8
XSTDFILL95_496 VDD VSS sg13g2_FILL8
XSTDFILL95_504 VDD VSS sg13g2_FILL8
XSTDFILL95_512 VDD VSS sg13g2_FILL8
XSTDFILL95_520 VDD VSS sg13g2_FILL8
XSTDFILL95_528 VDD VSS sg13g2_FILL8
XSTDFILL95_536 VDD VSS sg13g2_FILL8
XSTDFILL95_544 VDD VSS sg13g2_FILL8
XSTDFILL95_552 VDD VSS sg13g2_FILL8
XSTDFILL95_560 VDD VSS sg13g2_FILL8
XSTDFILL95_568 VDD VSS sg13g2_FILL8
XSTDFILL95_576 VDD VSS sg13g2_FILL8
XSTDFILL95_584 VDD VSS sg13g2_FILL8
XSTDFILL95_592 VDD VSS sg13g2_FILL8
XSTDFILL95_600 VDD VSS sg13g2_FILL8
XSTDFILL95_608 VDD VSS sg13g2_FILL8
XSTDFILL95_616 VDD VSS sg13g2_FILL8
XSTDFILL95_624 VDD VSS sg13g2_FILL8
XSTDFILL95_632 VDD VSS sg13g2_FILL8
XSTDFILL95_640 VDD VSS sg13g2_FILL8
XSTDFILL95_648 VDD VSS sg13g2_FILL8
XSTDFILL95_656 VDD VSS sg13g2_FILL8
XSTDFILL95_664 VDD VSS sg13g2_FILL8
XSTDFILL95_672 VDD VSS sg13g2_FILL8
XSTDFILL95_680 VDD VSS sg13g2_FILL8
XSTDFILL95_688 VDD VSS sg13g2_FILL8
XSTDFILL95_696 VDD VSS sg13g2_FILL8
XSTDFILL95_704 VDD VSS sg13g2_FILL8
XSTDFILL95_712 VDD VSS sg13g2_FILL8
XSTDFILL95_720 VDD VSS sg13g2_FILL8
XSTDFILL95_728 VDD VSS sg13g2_FILL8
XSTDFILL95_736 VDD VSS sg13g2_FILL8
XSTDFILL95_744 VDD VSS sg13g2_FILL8
XSTDFILL95_752 VDD VSS sg13g2_FILL8
XSTDFILL95_760 VDD VSS sg13g2_FILL8
XSTDFILL95_768 VDD VSS sg13g2_FILL8
XSTDFILL95_776 VDD VSS sg13g2_FILL8
XSTDFILL95_784 VDD VSS sg13g2_FILL8
XSTDFILL95_792 VDD VSS sg13g2_FILL8
XSTDFILL95_800 VDD VSS sg13g2_FILL8
XSTDFILL95_808 VDD VSS sg13g2_FILL8
XSTDFILL95_816 VDD VSS sg13g2_FILL8
XSTDFILL95_824 VDD VSS sg13g2_FILL8
XSTDFILL95_832 VDD VSS sg13g2_FILL8
XSTDFILL95_840 VDD VSS sg13g2_FILL8
XSTDFILL95_848 VDD VSS sg13g2_FILL8
XSTDFILL95_856 VDD VSS sg13g2_FILL8
XSTDFILL95_864 VDD VSS sg13g2_FILL8
XSTDFILL95_872 VDD VSS sg13g2_FILL8
XSTDFILL95_880 VDD VSS sg13g2_FILL8
XSTDFILL95_888 VDD VSS sg13g2_FILL8
XSTDFILL95_896 VDD VSS sg13g2_FILL8
XSTDFILL95_904 VDD VSS sg13g2_FILL8
XSTDFILL95_912 VDD VSS sg13g2_FILL8
XSTDFILL95_920 VDD VSS sg13g2_FILL8
XSTDFILL95_928 VDD VSS sg13g2_FILL8
XSTDFILL95_936 VDD VSS sg13g2_FILL8
XSTDFILL95_944 VDD VSS sg13g2_FILL8
XSTDFILL95_952 VDD VSS sg13g2_FILL8
XSTDFILL95_960 VDD VSS sg13g2_FILL8
XSTDFILL95_968 VDD VSS sg13g2_FILL8
XSTDFILL95_976 VDD VSS sg13g2_FILL8
XSTDFILL95_984 VDD VSS sg13g2_FILL8
XSTDFILL95_992 VDD VSS sg13g2_FILL8
XSTDFILL95_1000 VDD VSS sg13g2_FILL8
XSTDFILL95_1008 VDD VSS sg13g2_FILL8
XSTDFILL95_1016 VDD VSS sg13g2_FILL8
XSTDFILL95_1024 VDD VSS sg13g2_FILL8
XSTDFILL95_1032 VDD VSS sg13g2_FILL8
XSTDFILL95_1040 VDD VSS sg13g2_FILL8
XSTDFILL95_1048 VDD VSS sg13g2_FILL8
XSTDFILL95_1056 VDD VSS sg13g2_FILL8
XSTDFILL95_1064 VDD VSS sg13g2_FILL8
XSTDFILL95_1072 VDD VSS sg13g2_FILL8
XSTDFILL95_1080 VDD VSS sg13g2_FILL8
XSTDFILL95_1088 VDD VSS sg13g2_FILL8
XSTDFILL95_1096 VDD VSS sg13g2_FILL8
XSTDFILL95_1104 VDD VSS sg13g2_FILL8
XSTDFILL95_1112 VDD VSS sg13g2_FILL8
XSTDFILL95_1120 VDD VSS sg13g2_FILL8
XSTDFILL95_1128 VDD VSS sg13g2_FILL8
XSTDFILL95_1136 VDD VSS sg13g2_FILL8
XSTDFILL95_1144 VDD VSS sg13g2_FILL8
XSTDFILL95_1152 VDD VSS sg13g2_FILL8
XSTDFILL95_1160 VDD VSS sg13g2_FILL8
XSTDFILL95_1168 VDD VSS sg13g2_FILL8
XSTDFILL95_1176 VDD VSS sg13g2_FILL8
XSTDFILL95_1184 VDD VSS sg13g2_FILL8
XSTDFILL95_1192 VDD VSS sg13g2_FILL8
XSTDFILL95_1200 VDD VSS sg13g2_FILL8
XSTDFILL95_1208 VDD VSS sg13g2_FILL8
XSTDFILL95_1216 VDD VSS sg13g2_FILL8
XSTDFILL95_1224 VDD VSS sg13g2_FILL8
XSTDFILL95_1232 VDD VSS sg13g2_FILL8
XSTDFILL95_1240 VDD VSS sg13g2_FILL8
XSTDFILL95_1248 VDD VSS sg13g2_FILL8
XSTDFILL95_1256 VDD VSS sg13g2_FILL8
XSTDFILL95_1264 VDD VSS sg13g2_FILL8
XSTDFILL95_1272 VDD VSS sg13g2_FILL8
XSTDFILL95_1280 VDD VSS sg13g2_FILL8
XSTDFILL95_1288 VDD VSS sg13g2_FILL8
XSTDFILL95_1296 VDD VSS sg13g2_FILL8
XSTDFILL95_1304 VDD VSS sg13g2_FILL8
XSTDFILL95_1312 VDD VSS sg13g2_FILL8
XSTDFILL95_1320 VDD VSS sg13g2_FILL8
XSTDFILL95_1328 VDD VSS sg13g2_FILL8
XSTDFILL95_1336 VDD VSS sg13g2_FILL8
XSTDFILL95_1344 VDD VSS sg13g2_FILL8
XSTDFILL95_1352 VDD VSS sg13g2_FILL8
XSTDFILL95_1360 VDD VSS sg13g2_FILL8
XSTDFILL95_1368 VDD VSS sg13g2_FILL8
XSTDFILL95_1376 VDD VSS sg13g2_FILL8
XSTDFILL95_1384 VDD VSS sg13g2_FILL8
XSTDFILL95_1392 VDD VSS sg13g2_FILL8
XSTDFILL95_1400 VDD VSS sg13g2_FILL8
XSTDFILL95_1408 VDD VSS sg13g2_FILL8
XSTDFILL95_1416 VDD VSS sg13g2_FILL8
XSTDFILL95_1424 VDD VSS sg13g2_FILL8
XSTDFILL95_1432 VDD VSS sg13g2_FILL8
XSTDFILL95_1440 VDD VSS sg13g2_FILL8
XSTDFILL95_1448 VDD VSS sg13g2_FILL8
XSTDFILL95_1456 VDD VSS sg13g2_FILL8
XSTDFILL95_1464 VDD VSS sg13g2_FILL8
XSTDFILL95_1472 VDD VSS sg13g2_FILL8
XSTDFILL95_1480 VDD VSS sg13g2_FILL8
XSTDFILL95_1488 VDD VSS sg13g2_FILL8
XSTDFILL95_1496 VDD VSS sg13g2_FILL8
XSTDFILL95_1504 VDD VSS sg13g2_FILL8
XSTDFILL95_1512 VDD VSS sg13g2_FILL8
XSTDFILL95_1520 VDD VSS sg13g2_FILL8
XSTDFILL95_1528 VDD VSS sg13g2_FILL2
XSTDFILL95_1530 VDD VSS sg13g2_FILL1
XSTDFILL96_0 VDD VSS sg13g2_FILL8
XSTDFILL96_8 VDD VSS sg13g2_FILL8
XSTDFILL96_16 VDD VSS sg13g2_FILL8
XSTDFILL96_24 VDD VSS sg13g2_FILL8
XSTDFILL96_32 VDD VSS sg13g2_FILL8
XSTDFILL96_40 VDD VSS sg13g2_FILL8
XSTDFILL96_48 VDD VSS sg13g2_FILL8
XSTDFILL96_56 VDD VSS sg13g2_FILL8
XSTDFILL96_64 VDD VSS sg13g2_FILL8
XSTDFILL96_72 VDD VSS sg13g2_FILL8
XSTDFILL96_80 VDD VSS sg13g2_FILL8
XSTDFILL96_88 VDD VSS sg13g2_FILL8
XSTDFILL96_96 VDD VSS sg13g2_FILL8
XSTDFILL96_104 VDD VSS sg13g2_FILL8
XSTDFILL96_112 VDD VSS sg13g2_FILL8
XSTDFILL96_120 VDD VSS sg13g2_FILL8
XSTDFILL96_128 VDD VSS sg13g2_FILL8
XSTDFILL96_136 VDD VSS sg13g2_FILL8
XSTDFILL96_144 VDD VSS sg13g2_FILL8
XSTDFILL96_152 VDD VSS sg13g2_FILL8
XSTDFILL96_160 VDD VSS sg13g2_FILL8
XSTDFILL96_168 VDD VSS sg13g2_FILL8
XSTDFILL96_176 VDD VSS sg13g2_FILL8
XSTDFILL96_184 VDD VSS sg13g2_FILL8
XSTDFILL96_192 VDD VSS sg13g2_FILL8
XSTDFILL96_200 VDD VSS sg13g2_FILL8
XSTDFILL96_208 VDD VSS sg13g2_FILL8
XSTDFILL96_216 VDD VSS sg13g2_FILL8
XSTDFILL96_224 VDD VSS sg13g2_FILL8
XSTDFILL96_232 VDD VSS sg13g2_FILL8
XSTDFILL96_240 VDD VSS sg13g2_FILL8
XSTDFILL96_248 VDD VSS sg13g2_FILL8
XSTDFILL96_256 VDD VSS sg13g2_FILL8
XSTDFILL96_264 VDD VSS sg13g2_FILL8
XSTDFILL96_272 VDD VSS sg13g2_FILL8
XSTDFILL96_280 VDD VSS sg13g2_FILL8
XSTDFILL96_288 VDD VSS sg13g2_FILL8
XSTDFILL96_296 VDD VSS sg13g2_FILL8
XSTDFILL96_304 VDD VSS sg13g2_FILL8
XSTDFILL96_312 VDD VSS sg13g2_FILL8
XSTDFILL96_320 VDD VSS sg13g2_FILL8
XSTDFILL96_328 VDD VSS sg13g2_FILL8
XSTDFILL96_336 VDD VSS sg13g2_FILL8
XSTDFILL96_344 VDD VSS sg13g2_FILL8
XSTDFILL96_352 VDD VSS sg13g2_FILL8
XSTDFILL96_360 VDD VSS sg13g2_FILL8
XSTDFILL96_368 VDD VSS sg13g2_FILL8
XSTDFILL96_376 VDD VSS sg13g2_FILL8
XSTDFILL96_384 VDD VSS sg13g2_FILL8
XSTDFILL96_392 VDD VSS sg13g2_FILL8
XSTDFILL96_400 VDD VSS sg13g2_FILL8
XSTDFILL96_408 VDD VSS sg13g2_FILL8
XSTDFILL96_416 VDD VSS sg13g2_FILL8
XSTDFILL96_424 VDD VSS sg13g2_FILL8
XSTDFILL96_432 VDD VSS sg13g2_FILL8
XSTDFILL96_440 VDD VSS sg13g2_FILL8
XSTDFILL96_448 VDD VSS sg13g2_FILL8
XSTDFILL96_456 VDD VSS sg13g2_FILL8
XSTDFILL96_464 VDD VSS sg13g2_FILL8
XSTDFILL96_472 VDD VSS sg13g2_FILL8
XSTDFILL96_480 VDD VSS sg13g2_FILL8
XSTDFILL96_488 VDD VSS sg13g2_FILL8
XSTDFILL96_496 VDD VSS sg13g2_FILL8
XSTDFILL96_504 VDD VSS sg13g2_FILL8
XSTDFILL96_512 VDD VSS sg13g2_FILL8
XSTDFILL96_520 VDD VSS sg13g2_FILL8
XSTDFILL96_528 VDD VSS sg13g2_FILL8
XSTDFILL96_536 VDD VSS sg13g2_FILL8
XSTDFILL96_544 VDD VSS sg13g2_FILL8
XSTDFILL96_552 VDD VSS sg13g2_FILL8
XSTDFILL96_560 VDD VSS sg13g2_FILL8
XSTDFILL96_568 VDD VSS sg13g2_FILL8
XSTDFILL96_576 VDD VSS sg13g2_FILL8
XSTDFILL96_584 VDD VSS sg13g2_FILL8
XSTDFILL96_592 VDD VSS sg13g2_FILL8
XSTDFILL96_600 VDD VSS sg13g2_FILL8
XSTDFILL96_608 VDD VSS sg13g2_FILL8
XSTDFILL96_616 VDD VSS sg13g2_FILL8
XSTDFILL96_624 VDD VSS sg13g2_FILL8
XSTDFILL96_632 VDD VSS sg13g2_FILL8
XSTDFILL96_640 VDD VSS sg13g2_FILL8
XSTDFILL96_648 VDD VSS sg13g2_FILL8
XSTDFILL96_656 VDD VSS sg13g2_FILL8
XSTDFILL96_664 VDD VSS sg13g2_FILL8
XSTDFILL96_672 VDD VSS sg13g2_FILL8
XSTDFILL96_680 VDD VSS sg13g2_FILL8
XSTDFILL96_688 VDD VSS sg13g2_FILL8
XSTDFILL96_696 VDD VSS sg13g2_FILL8
XSTDFILL96_704 VDD VSS sg13g2_FILL8
XSTDFILL96_712 VDD VSS sg13g2_FILL8
XSTDFILL96_720 VDD VSS sg13g2_FILL8
XSTDFILL96_728 VDD VSS sg13g2_FILL8
XSTDFILL96_736 VDD VSS sg13g2_FILL8
XSTDFILL96_744 VDD VSS sg13g2_FILL8
XSTDFILL96_752 VDD VSS sg13g2_FILL8
XSTDFILL96_760 VDD VSS sg13g2_FILL8
XSTDFILL96_768 VDD VSS sg13g2_FILL8
XSTDFILL96_776 VDD VSS sg13g2_FILL8
XSTDFILL96_784 VDD VSS sg13g2_FILL8
XSTDFILL96_792 VDD VSS sg13g2_FILL8
XSTDFILL96_800 VDD VSS sg13g2_FILL8
XSTDFILL96_808 VDD VSS sg13g2_FILL8
XSTDFILL96_816 VDD VSS sg13g2_FILL8
XSTDFILL96_824 VDD VSS sg13g2_FILL8
XSTDFILL96_832 VDD VSS sg13g2_FILL8
XSTDFILL96_840 VDD VSS sg13g2_FILL8
XSTDFILL96_848 VDD VSS sg13g2_FILL8
XSTDFILL96_856 VDD VSS sg13g2_FILL8
XSTDFILL96_864 VDD VSS sg13g2_FILL8
XSTDFILL96_872 VDD VSS sg13g2_FILL8
XSTDFILL96_880 VDD VSS sg13g2_FILL8
XSTDFILL96_888 VDD VSS sg13g2_FILL8
XSTDFILL96_896 VDD VSS sg13g2_FILL8
XSTDFILL96_904 VDD VSS sg13g2_FILL8
XSTDFILL96_912 VDD VSS sg13g2_FILL8
XSTDFILL96_920 VDD VSS sg13g2_FILL8
XSTDFILL96_928 VDD VSS sg13g2_FILL8
XSTDFILL96_936 VDD VSS sg13g2_FILL8
XSTDFILL96_944 VDD VSS sg13g2_FILL8
XSTDFILL96_952 VDD VSS sg13g2_FILL8
XSTDFILL96_960 VDD VSS sg13g2_FILL8
XSTDFILL96_968 VDD VSS sg13g2_FILL8
XSTDFILL96_976 VDD VSS sg13g2_FILL8
XSTDFILL96_984 VDD VSS sg13g2_FILL8
XSTDFILL96_992 VDD VSS sg13g2_FILL8
XSTDFILL96_1000 VDD VSS sg13g2_FILL8
XSTDFILL96_1008 VDD VSS sg13g2_FILL8
XSTDFILL96_1016 VDD VSS sg13g2_FILL8
XSTDFILL96_1024 VDD VSS sg13g2_FILL8
XSTDFILL96_1032 VDD VSS sg13g2_FILL8
XSTDFILL96_1040 VDD VSS sg13g2_FILL8
XSTDFILL96_1048 VDD VSS sg13g2_FILL8
XSTDFILL96_1056 VDD VSS sg13g2_FILL8
XSTDFILL96_1064 VDD VSS sg13g2_FILL8
XSTDFILL96_1072 VDD VSS sg13g2_FILL8
XSTDFILL96_1080 VDD VSS sg13g2_FILL8
XSTDFILL96_1088 VDD VSS sg13g2_FILL8
XSTDFILL96_1096 VDD VSS sg13g2_FILL8
XSTDFILL96_1104 VDD VSS sg13g2_FILL8
XSTDFILL96_1112 VDD VSS sg13g2_FILL8
XSTDFILL96_1120 VDD VSS sg13g2_FILL8
XSTDFILL96_1128 VDD VSS sg13g2_FILL8
XSTDFILL96_1136 VDD VSS sg13g2_FILL8
XSTDFILL96_1144 VDD VSS sg13g2_FILL8
XSTDFILL96_1152 VDD VSS sg13g2_FILL8
XSTDFILL96_1160 VDD VSS sg13g2_FILL8
XSTDFILL96_1168 VDD VSS sg13g2_FILL8
XSTDFILL96_1176 VDD VSS sg13g2_FILL8
XSTDFILL96_1184 VDD VSS sg13g2_FILL8
XSTDFILL96_1192 VDD VSS sg13g2_FILL8
XSTDFILL96_1200 VDD VSS sg13g2_FILL8
XSTDFILL96_1208 VDD VSS sg13g2_FILL8
XSTDFILL96_1216 VDD VSS sg13g2_FILL8
XSTDFILL96_1224 VDD VSS sg13g2_FILL8
XSTDFILL96_1232 VDD VSS sg13g2_FILL8
XSTDFILL96_1240 VDD VSS sg13g2_FILL8
XSTDFILL96_1248 VDD VSS sg13g2_FILL8
XSTDFILL96_1256 VDD VSS sg13g2_FILL8
XSTDFILL96_1264 VDD VSS sg13g2_FILL8
XSTDFILL96_1272 VDD VSS sg13g2_FILL8
XSTDFILL96_1280 VDD VSS sg13g2_FILL8
XSTDFILL96_1288 VDD VSS sg13g2_FILL8
XSTDFILL96_1296 VDD VSS sg13g2_FILL8
XSTDFILL96_1304 VDD VSS sg13g2_FILL8
XSTDFILL96_1312 VDD VSS sg13g2_FILL8
XSTDFILL96_1320 VDD VSS sg13g2_FILL8
XSTDFILL96_1328 VDD VSS sg13g2_FILL8
XSTDFILL96_1336 VDD VSS sg13g2_FILL8
XSTDFILL96_1344 VDD VSS sg13g2_FILL8
XSTDFILL96_1352 VDD VSS sg13g2_FILL8
XSTDFILL96_1360 VDD VSS sg13g2_FILL8
XSTDFILL96_1368 VDD VSS sg13g2_FILL8
XSTDFILL96_1376 VDD VSS sg13g2_FILL8
XSTDFILL96_1384 VDD VSS sg13g2_FILL8
XSTDFILL96_1392 VDD VSS sg13g2_FILL8
XSTDFILL96_1400 VDD VSS sg13g2_FILL8
XSTDFILL96_1408 VDD VSS sg13g2_FILL8
XSTDFILL96_1416 VDD VSS sg13g2_FILL8
XSTDFILL96_1424 VDD VSS sg13g2_FILL8
XSTDFILL96_1432 VDD VSS sg13g2_FILL8
XSTDFILL96_1440 VDD VSS sg13g2_FILL8
XSTDFILL96_1448 VDD VSS sg13g2_FILL8
XSTDFILL96_1456 VDD VSS sg13g2_FILL8
XSTDFILL96_1464 VDD VSS sg13g2_FILL8
XSTDFILL96_1472 VDD VSS sg13g2_FILL8
XSTDFILL96_1480 VDD VSS sg13g2_FILL8
XSTDFILL96_1488 VDD VSS sg13g2_FILL8
XSTDFILL96_1496 VDD VSS sg13g2_FILL8
XSTDFILL96_1504 VDD VSS sg13g2_FILL8
XSTDFILL96_1512 VDD VSS sg13g2_FILL8
XSTDFILL96_1520 VDD VSS sg13g2_FILL8
XSTDFILL96_1528 VDD VSS sg13g2_FILL2
XSTDFILL96_1530 VDD VSS sg13g2_FILL1
XSTDFILL97_0 VDD VSS sg13g2_FILL8
XSTDFILL97_8 VDD VSS sg13g2_FILL8
XSTDFILL97_16 VDD VSS sg13g2_FILL8
XSTDFILL97_24 VDD VSS sg13g2_FILL8
XSTDFILL97_32 VDD VSS sg13g2_FILL8
XSTDFILL97_40 VDD VSS sg13g2_FILL8
XSTDFILL97_48 VDD VSS sg13g2_FILL8
XSTDFILL97_56 VDD VSS sg13g2_FILL8
XSTDFILL97_64 VDD VSS sg13g2_FILL8
XSTDFILL97_72 VDD VSS sg13g2_FILL8
XSTDFILL97_80 VDD VSS sg13g2_FILL8
XSTDFILL97_88 VDD VSS sg13g2_FILL8
XSTDFILL97_96 VDD VSS sg13g2_FILL8
XSTDFILL97_104 VDD VSS sg13g2_FILL8
XSTDFILL97_112 VDD VSS sg13g2_FILL8
XSTDFILL97_120 VDD VSS sg13g2_FILL8
XSTDFILL97_128 VDD VSS sg13g2_FILL8
XSTDFILL97_136 VDD VSS sg13g2_FILL8
XSTDFILL97_144 VDD VSS sg13g2_FILL8
XSTDFILL97_152 VDD VSS sg13g2_FILL8
XSTDFILL97_160 VDD VSS sg13g2_FILL8
XSTDFILL97_168 VDD VSS sg13g2_FILL8
XSTDFILL97_176 VDD VSS sg13g2_FILL8
XSTDFILL97_184 VDD VSS sg13g2_FILL8
XSTDFILL97_192 VDD VSS sg13g2_FILL8
XSTDFILL97_200 VDD VSS sg13g2_FILL8
XSTDFILL97_208 VDD VSS sg13g2_FILL8
XSTDFILL97_216 VDD VSS sg13g2_FILL8
XSTDFILL97_224 VDD VSS sg13g2_FILL8
XSTDFILL97_232 VDD VSS sg13g2_FILL8
XSTDFILL97_240 VDD VSS sg13g2_FILL8
XSTDFILL97_248 VDD VSS sg13g2_FILL8
XSTDFILL97_256 VDD VSS sg13g2_FILL8
XSTDFILL97_264 VDD VSS sg13g2_FILL8
XSTDFILL97_272 VDD VSS sg13g2_FILL8
XSTDFILL97_280 VDD VSS sg13g2_FILL8
XSTDFILL97_288 VDD VSS sg13g2_FILL8
XSTDFILL97_296 VDD VSS sg13g2_FILL8
XSTDFILL97_304 VDD VSS sg13g2_FILL8
XSTDFILL97_312 VDD VSS sg13g2_FILL8
XSTDFILL97_320 VDD VSS sg13g2_FILL8
XSTDFILL97_328 VDD VSS sg13g2_FILL8
XSTDFILL97_336 VDD VSS sg13g2_FILL8
XSTDFILL97_344 VDD VSS sg13g2_FILL8
XSTDFILL97_352 VDD VSS sg13g2_FILL8
XSTDFILL97_360 VDD VSS sg13g2_FILL8
XSTDFILL97_368 VDD VSS sg13g2_FILL8
XSTDFILL97_376 VDD VSS sg13g2_FILL8
XSTDFILL97_384 VDD VSS sg13g2_FILL8
XSTDFILL97_392 VDD VSS sg13g2_FILL8
XSTDFILL97_400 VDD VSS sg13g2_FILL8
XSTDFILL97_408 VDD VSS sg13g2_FILL8
XSTDFILL97_416 VDD VSS sg13g2_FILL8
XSTDFILL97_424 VDD VSS sg13g2_FILL8
XSTDFILL97_432 VDD VSS sg13g2_FILL8
XSTDFILL97_440 VDD VSS sg13g2_FILL8
XSTDFILL97_448 VDD VSS sg13g2_FILL8
XSTDFILL97_456 VDD VSS sg13g2_FILL8
XSTDFILL97_464 VDD VSS sg13g2_FILL8
XSTDFILL97_472 VDD VSS sg13g2_FILL8
XSTDFILL97_480 VDD VSS sg13g2_FILL8
XSTDFILL97_488 VDD VSS sg13g2_FILL8
XSTDFILL97_496 VDD VSS sg13g2_FILL8
XSTDFILL97_504 VDD VSS sg13g2_FILL8
XSTDFILL97_512 VDD VSS sg13g2_FILL8
XSTDFILL97_520 VDD VSS sg13g2_FILL8
XSTDFILL97_528 VDD VSS sg13g2_FILL8
XSTDFILL97_536 VDD VSS sg13g2_FILL8
XSTDFILL97_544 VDD VSS sg13g2_FILL8
XSTDFILL97_552 VDD VSS sg13g2_FILL8
XSTDFILL97_560 VDD VSS sg13g2_FILL8
XSTDFILL97_568 VDD VSS sg13g2_FILL8
XSTDFILL97_576 VDD VSS sg13g2_FILL8
XSTDFILL97_584 VDD VSS sg13g2_FILL8
XSTDFILL97_592 VDD VSS sg13g2_FILL8
XSTDFILL97_600 VDD VSS sg13g2_FILL8
XSTDFILL97_608 VDD VSS sg13g2_FILL8
XSTDFILL97_616 VDD VSS sg13g2_FILL8
XSTDFILL97_624 VDD VSS sg13g2_FILL8
XSTDFILL97_632 VDD VSS sg13g2_FILL8
XSTDFILL97_640 VDD VSS sg13g2_FILL8
XSTDFILL97_648 VDD VSS sg13g2_FILL8
XSTDFILL97_656 VDD VSS sg13g2_FILL8
XSTDFILL97_664 VDD VSS sg13g2_FILL8
XSTDFILL97_672 VDD VSS sg13g2_FILL8
XSTDFILL97_680 VDD VSS sg13g2_FILL8
XSTDFILL97_688 VDD VSS sg13g2_FILL8
XSTDFILL97_696 VDD VSS sg13g2_FILL8
XSTDFILL97_704 VDD VSS sg13g2_FILL8
XSTDFILL97_712 VDD VSS sg13g2_FILL8
XSTDFILL97_720 VDD VSS sg13g2_FILL8
XSTDFILL97_728 VDD VSS sg13g2_FILL8
XSTDFILL97_736 VDD VSS sg13g2_FILL8
XSTDFILL97_744 VDD VSS sg13g2_FILL8
XSTDFILL97_752 VDD VSS sg13g2_FILL8
XSTDFILL97_760 VDD VSS sg13g2_FILL8
XSTDFILL97_768 VDD VSS sg13g2_FILL8
XSTDFILL97_776 VDD VSS sg13g2_FILL8
XSTDFILL97_784 VDD VSS sg13g2_FILL8
XSTDFILL97_792 VDD VSS sg13g2_FILL8
XSTDFILL97_800 VDD VSS sg13g2_FILL8
XSTDFILL97_808 VDD VSS sg13g2_FILL8
XSTDFILL97_816 VDD VSS sg13g2_FILL8
XSTDFILL97_824 VDD VSS sg13g2_FILL8
XSTDFILL97_832 VDD VSS sg13g2_FILL8
XSTDFILL97_840 VDD VSS sg13g2_FILL8
XSTDFILL97_848 VDD VSS sg13g2_FILL8
XSTDFILL97_856 VDD VSS sg13g2_FILL8
XSTDFILL97_864 VDD VSS sg13g2_FILL8
XSTDFILL97_872 VDD VSS sg13g2_FILL8
XSTDFILL97_880 VDD VSS sg13g2_FILL8
XSTDFILL97_888 VDD VSS sg13g2_FILL8
XSTDFILL97_896 VDD VSS sg13g2_FILL8
XSTDFILL97_904 VDD VSS sg13g2_FILL8
XSTDFILL97_912 VDD VSS sg13g2_FILL8
XSTDFILL97_920 VDD VSS sg13g2_FILL8
XSTDFILL97_928 VDD VSS sg13g2_FILL8
XSTDFILL97_936 VDD VSS sg13g2_FILL8
XSTDFILL97_944 VDD VSS sg13g2_FILL8
XSTDFILL97_952 VDD VSS sg13g2_FILL8
XSTDFILL97_960 VDD VSS sg13g2_FILL8
XSTDFILL97_968 VDD VSS sg13g2_FILL8
XSTDFILL97_976 VDD VSS sg13g2_FILL8
XSTDFILL97_984 VDD VSS sg13g2_FILL8
XSTDFILL97_992 VDD VSS sg13g2_FILL8
XSTDFILL97_1000 VDD VSS sg13g2_FILL8
XSTDFILL97_1008 VDD VSS sg13g2_FILL8
XSTDFILL97_1016 VDD VSS sg13g2_FILL8
XSTDFILL97_1024 VDD VSS sg13g2_FILL8
XSTDFILL97_1032 VDD VSS sg13g2_FILL8
XSTDFILL97_1040 VDD VSS sg13g2_FILL8
XSTDFILL97_1048 VDD VSS sg13g2_FILL8
XSTDFILL97_1056 VDD VSS sg13g2_FILL8
XSTDFILL97_1064 VDD VSS sg13g2_FILL8
XSTDFILL97_1072 VDD VSS sg13g2_FILL8
XSTDFILL97_1080 VDD VSS sg13g2_FILL8
XSTDFILL97_1088 VDD VSS sg13g2_FILL8
XSTDFILL97_1096 VDD VSS sg13g2_FILL8
XSTDFILL97_1104 VDD VSS sg13g2_FILL8
XSTDFILL97_1112 VDD VSS sg13g2_FILL8
XSTDFILL97_1120 VDD VSS sg13g2_FILL8
XSTDFILL97_1128 VDD VSS sg13g2_FILL8
XSTDFILL97_1136 VDD VSS sg13g2_FILL8
XSTDFILL97_1144 VDD VSS sg13g2_FILL8
XSTDFILL97_1152 VDD VSS sg13g2_FILL8
XSTDFILL97_1160 VDD VSS sg13g2_FILL8
XSTDFILL97_1168 VDD VSS sg13g2_FILL8
XSTDFILL97_1176 VDD VSS sg13g2_FILL8
XSTDFILL97_1184 VDD VSS sg13g2_FILL8
XSTDFILL97_1192 VDD VSS sg13g2_FILL8
XSTDFILL97_1200 VDD VSS sg13g2_FILL8
XSTDFILL97_1208 VDD VSS sg13g2_FILL8
XSTDFILL97_1216 VDD VSS sg13g2_FILL8
XSTDFILL97_1224 VDD VSS sg13g2_FILL8
XSTDFILL97_1232 VDD VSS sg13g2_FILL8
XSTDFILL97_1240 VDD VSS sg13g2_FILL8
XSTDFILL97_1248 VDD VSS sg13g2_FILL8
XSTDFILL97_1256 VDD VSS sg13g2_FILL8
XSTDFILL97_1264 VDD VSS sg13g2_FILL8
XSTDFILL97_1272 VDD VSS sg13g2_FILL8
XSTDFILL97_1280 VDD VSS sg13g2_FILL8
XSTDFILL97_1288 VDD VSS sg13g2_FILL8
XSTDFILL97_1296 VDD VSS sg13g2_FILL8
XSTDFILL97_1304 VDD VSS sg13g2_FILL8
XSTDFILL97_1312 VDD VSS sg13g2_FILL8
XSTDFILL97_1320 VDD VSS sg13g2_FILL8
XSTDFILL97_1328 VDD VSS sg13g2_FILL8
XSTDFILL97_1336 VDD VSS sg13g2_FILL8
XSTDFILL97_1344 VDD VSS sg13g2_FILL8
XSTDFILL97_1352 VDD VSS sg13g2_FILL8
XSTDFILL97_1360 VDD VSS sg13g2_FILL8
XSTDFILL97_1368 VDD VSS sg13g2_FILL8
XSTDFILL97_1376 VDD VSS sg13g2_FILL8
XSTDFILL97_1384 VDD VSS sg13g2_FILL8
XSTDFILL97_1392 VDD VSS sg13g2_FILL8
XSTDFILL97_1400 VDD VSS sg13g2_FILL8
XSTDFILL97_1408 VDD VSS sg13g2_FILL8
XSTDFILL97_1416 VDD VSS sg13g2_FILL8
XSTDFILL97_1424 VDD VSS sg13g2_FILL8
XSTDFILL97_1432 VDD VSS sg13g2_FILL8
XSTDFILL97_1440 VDD VSS sg13g2_FILL8
XSTDFILL97_1448 VDD VSS sg13g2_FILL8
XSTDFILL97_1456 VDD VSS sg13g2_FILL8
XSTDFILL97_1464 VDD VSS sg13g2_FILL8
XSTDFILL97_1472 VDD VSS sg13g2_FILL8
XSTDFILL97_1480 VDD VSS sg13g2_FILL8
XSTDFILL97_1488 VDD VSS sg13g2_FILL8
XSTDFILL97_1496 VDD VSS sg13g2_FILL8
XSTDFILL97_1504 VDD VSS sg13g2_FILL8
XSTDFILL97_1512 VDD VSS sg13g2_FILL8
XSTDFILL97_1520 VDD VSS sg13g2_FILL8
XSTDFILL97_1528 VDD VSS sg13g2_FILL2
XSTDFILL97_1530 VDD VSS sg13g2_FILL1
XSTDFILL98_0 VDD VSS sg13g2_FILL8
XSTDFILL98_8 VDD VSS sg13g2_FILL8
XSTDFILL98_16 VDD VSS sg13g2_FILL8
XSTDFILL98_24 VDD VSS sg13g2_FILL8
XSTDFILL98_32 VDD VSS sg13g2_FILL8
XSTDFILL98_40 VDD VSS sg13g2_FILL8
XSTDFILL98_48 VDD VSS sg13g2_FILL8
XSTDFILL98_56 VDD VSS sg13g2_FILL8
XSTDFILL98_64 VDD VSS sg13g2_FILL8
XSTDFILL98_72 VDD VSS sg13g2_FILL8
XSTDFILL98_80 VDD VSS sg13g2_FILL8
XSTDFILL98_88 VDD VSS sg13g2_FILL8
XSTDFILL98_96 VDD VSS sg13g2_FILL8
XSTDFILL98_104 VDD VSS sg13g2_FILL8
XSTDFILL98_112 VDD VSS sg13g2_FILL8
XSTDFILL98_120 VDD VSS sg13g2_FILL8
XSTDFILL98_128 VDD VSS sg13g2_FILL8
XSTDFILL98_136 VDD VSS sg13g2_FILL8
XSTDFILL98_144 VDD VSS sg13g2_FILL8
XSTDFILL98_152 VDD VSS sg13g2_FILL8
XSTDFILL98_160 VDD VSS sg13g2_FILL8
XSTDFILL98_168 VDD VSS sg13g2_FILL8
XSTDFILL98_176 VDD VSS sg13g2_FILL8
XSTDFILL98_184 VDD VSS sg13g2_FILL8
XSTDFILL98_192 VDD VSS sg13g2_FILL8
XSTDFILL98_200 VDD VSS sg13g2_FILL8
XSTDFILL98_208 VDD VSS sg13g2_FILL8
XSTDFILL98_216 VDD VSS sg13g2_FILL8
XSTDFILL98_224 VDD VSS sg13g2_FILL8
XSTDFILL98_232 VDD VSS sg13g2_FILL8
XSTDFILL98_240 VDD VSS sg13g2_FILL8
XSTDFILL98_248 VDD VSS sg13g2_FILL8
XSTDFILL98_256 VDD VSS sg13g2_FILL8
XSTDFILL98_264 VDD VSS sg13g2_FILL8
XSTDFILL98_272 VDD VSS sg13g2_FILL8
XSTDFILL98_280 VDD VSS sg13g2_FILL8
XSTDFILL98_288 VDD VSS sg13g2_FILL8
XSTDFILL98_296 VDD VSS sg13g2_FILL8
XSTDFILL98_304 VDD VSS sg13g2_FILL8
XSTDFILL98_312 VDD VSS sg13g2_FILL8
XSTDFILL98_320 VDD VSS sg13g2_FILL8
XSTDFILL98_328 VDD VSS sg13g2_FILL8
XSTDFILL98_336 VDD VSS sg13g2_FILL8
XSTDFILL98_344 VDD VSS sg13g2_FILL8
XSTDFILL98_352 VDD VSS sg13g2_FILL8
XSTDFILL98_360 VDD VSS sg13g2_FILL8
XSTDFILL98_368 VDD VSS sg13g2_FILL8
XSTDFILL98_376 VDD VSS sg13g2_FILL8
XSTDFILL98_384 VDD VSS sg13g2_FILL8
XSTDFILL98_392 VDD VSS sg13g2_FILL8
XSTDFILL98_400 VDD VSS sg13g2_FILL8
XSTDFILL98_408 VDD VSS sg13g2_FILL8
XSTDFILL98_416 VDD VSS sg13g2_FILL8
XSTDFILL98_424 VDD VSS sg13g2_FILL8
XSTDFILL98_432 VDD VSS sg13g2_FILL8
XSTDFILL98_440 VDD VSS sg13g2_FILL8
XSTDFILL98_448 VDD VSS sg13g2_FILL8
XSTDFILL98_456 VDD VSS sg13g2_FILL8
XSTDFILL98_464 VDD VSS sg13g2_FILL8
XSTDFILL98_472 VDD VSS sg13g2_FILL8
XSTDFILL98_480 VDD VSS sg13g2_FILL8
XSTDFILL98_488 VDD VSS sg13g2_FILL8
XSTDFILL98_496 VDD VSS sg13g2_FILL8
XSTDFILL98_504 VDD VSS sg13g2_FILL8
XSTDFILL98_512 VDD VSS sg13g2_FILL8
XSTDFILL98_520 VDD VSS sg13g2_FILL8
XSTDFILL98_528 VDD VSS sg13g2_FILL8
XSTDFILL98_536 VDD VSS sg13g2_FILL8
XSTDFILL98_544 VDD VSS sg13g2_FILL8
XSTDFILL98_552 VDD VSS sg13g2_FILL8
XSTDFILL98_560 VDD VSS sg13g2_FILL8
XSTDFILL98_568 VDD VSS sg13g2_FILL8
XSTDFILL98_576 VDD VSS sg13g2_FILL8
XSTDFILL98_584 VDD VSS sg13g2_FILL8
XSTDFILL98_592 VDD VSS sg13g2_FILL8
XSTDFILL98_600 VDD VSS sg13g2_FILL8
XSTDFILL98_608 VDD VSS sg13g2_FILL8
XSTDFILL98_616 VDD VSS sg13g2_FILL8
XSTDFILL98_624 VDD VSS sg13g2_FILL8
XSTDFILL98_632 VDD VSS sg13g2_FILL8
XSTDFILL98_640 VDD VSS sg13g2_FILL8
XSTDFILL98_648 VDD VSS sg13g2_FILL8
XSTDFILL98_656 VDD VSS sg13g2_FILL8
XSTDFILL98_664 VDD VSS sg13g2_FILL8
XSTDFILL98_672 VDD VSS sg13g2_FILL8
XSTDFILL98_680 VDD VSS sg13g2_FILL8
XSTDFILL98_688 VDD VSS sg13g2_FILL8
XSTDFILL98_696 VDD VSS sg13g2_FILL8
XSTDFILL98_704 VDD VSS sg13g2_FILL8
XSTDFILL98_712 VDD VSS sg13g2_FILL8
XSTDFILL98_720 VDD VSS sg13g2_FILL8
XSTDFILL98_728 VDD VSS sg13g2_FILL8
XSTDFILL98_736 VDD VSS sg13g2_FILL8
XSTDFILL98_744 VDD VSS sg13g2_FILL8
XSTDFILL98_752 VDD VSS sg13g2_FILL8
XSTDFILL98_760 VDD VSS sg13g2_FILL8
XSTDFILL98_768 VDD VSS sg13g2_FILL8
XSTDFILL98_776 VDD VSS sg13g2_FILL8
XSTDFILL98_784 VDD VSS sg13g2_FILL8
XSTDFILL98_792 VDD VSS sg13g2_FILL8
XSTDFILL98_800 VDD VSS sg13g2_FILL8
XSTDFILL98_808 VDD VSS sg13g2_FILL8
XSTDFILL98_816 VDD VSS sg13g2_FILL8
XSTDFILL98_824 VDD VSS sg13g2_FILL8
XSTDFILL98_832 VDD VSS sg13g2_FILL8
XSTDFILL98_840 VDD VSS sg13g2_FILL8
XSTDFILL98_848 VDD VSS sg13g2_FILL8
XSTDFILL98_856 VDD VSS sg13g2_FILL8
XSTDFILL98_864 VDD VSS sg13g2_FILL8
XSTDFILL98_872 VDD VSS sg13g2_FILL8
XSTDFILL98_880 VDD VSS sg13g2_FILL8
XSTDFILL98_888 VDD VSS sg13g2_FILL8
XSTDFILL98_896 VDD VSS sg13g2_FILL8
XSTDFILL98_904 VDD VSS sg13g2_FILL8
XSTDFILL98_912 VDD VSS sg13g2_FILL8
XSTDFILL98_920 VDD VSS sg13g2_FILL8
XSTDFILL98_928 VDD VSS sg13g2_FILL8
XSTDFILL98_936 VDD VSS sg13g2_FILL8
XSTDFILL98_944 VDD VSS sg13g2_FILL8
XSTDFILL98_952 VDD VSS sg13g2_FILL8
XSTDFILL98_960 VDD VSS sg13g2_FILL8
XSTDFILL98_968 VDD VSS sg13g2_FILL8
XSTDFILL98_976 VDD VSS sg13g2_FILL8
XSTDFILL98_984 VDD VSS sg13g2_FILL8
XSTDFILL98_992 VDD VSS sg13g2_FILL8
XSTDFILL98_1000 VDD VSS sg13g2_FILL8
XSTDFILL98_1008 VDD VSS sg13g2_FILL8
XSTDFILL98_1016 VDD VSS sg13g2_FILL8
XSTDFILL98_1024 VDD VSS sg13g2_FILL8
XSTDFILL98_1032 VDD VSS sg13g2_FILL8
XSTDFILL98_1040 VDD VSS sg13g2_FILL8
XSTDFILL98_1048 VDD VSS sg13g2_FILL8
XSTDFILL98_1056 VDD VSS sg13g2_FILL8
XSTDFILL98_1064 VDD VSS sg13g2_FILL8
XSTDFILL98_1072 VDD VSS sg13g2_FILL8
XSTDFILL98_1080 VDD VSS sg13g2_FILL8
XSTDFILL98_1088 VDD VSS sg13g2_FILL8
XSTDFILL98_1096 VDD VSS sg13g2_FILL8
XSTDFILL98_1104 VDD VSS sg13g2_FILL8
XSTDFILL98_1112 VDD VSS sg13g2_FILL8
XSTDFILL98_1120 VDD VSS sg13g2_FILL8
XSTDFILL98_1128 VDD VSS sg13g2_FILL8
XSTDFILL98_1136 VDD VSS sg13g2_FILL8
XSTDFILL98_1144 VDD VSS sg13g2_FILL8
XSTDFILL98_1152 VDD VSS sg13g2_FILL8
XSTDFILL98_1160 VDD VSS sg13g2_FILL8
XSTDFILL98_1168 VDD VSS sg13g2_FILL8
XSTDFILL98_1176 VDD VSS sg13g2_FILL8
XSTDFILL98_1184 VDD VSS sg13g2_FILL8
XSTDFILL98_1192 VDD VSS sg13g2_FILL8
XSTDFILL98_1200 VDD VSS sg13g2_FILL8
XSTDFILL98_1208 VDD VSS sg13g2_FILL8
XSTDFILL98_1216 VDD VSS sg13g2_FILL8
XSTDFILL98_1224 VDD VSS sg13g2_FILL8
XSTDFILL98_1232 VDD VSS sg13g2_FILL8
XSTDFILL98_1240 VDD VSS sg13g2_FILL8
XSTDFILL98_1248 VDD VSS sg13g2_FILL8
XSTDFILL98_1256 VDD VSS sg13g2_FILL8
XSTDFILL98_1264 VDD VSS sg13g2_FILL8
XSTDFILL98_1272 VDD VSS sg13g2_FILL8
XSTDFILL98_1280 VDD VSS sg13g2_FILL8
XSTDFILL98_1288 VDD VSS sg13g2_FILL8
XSTDFILL98_1296 VDD VSS sg13g2_FILL8
XSTDFILL98_1304 VDD VSS sg13g2_FILL8
XSTDFILL98_1312 VDD VSS sg13g2_FILL8
XSTDFILL98_1320 VDD VSS sg13g2_FILL8
XSTDFILL98_1328 VDD VSS sg13g2_FILL8
XSTDFILL98_1336 VDD VSS sg13g2_FILL8
XSTDFILL98_1344 VDD VSS sg13g2_FILL8
XSTDFILL98_1352 VDD VSS sg13g2_FILL8
XSTDFILL98_1360 VDD VSS sg13g2_FILL8
XSTDFILL98_1368 VDD VSS sg13g2_FILL8
XSTDFILL98_1376 VDD VSS sg13g2_FILL8
XSTDFILL98_1384 VDD VSS sg13g2_FILL8
XSTDFILL98_1392 VDD VSS sg13g2_FILL8
XSTDFILL98_1400 VDD VSS sg13g2_FILL8
XSTDFILL98_1408 VDD VSS sg13g2_FILL8
XSTDFILL98_1416 VDD VSS sg13g2_FILL8
XSTDFILL98_1424 VDD VSS sg13g2_FILL8
XSTDFILL98_1432 VDD VSS sg13g2_FILL8
XSTDFILL98_1440 VDD VSS sg13g2_FILL8
XSTDFILL98_1448 VDD VSS sg13g2_FILL8
XSTDFILL98_1456 VDD VSS sg13g2_FILL8
XSTDFILL98_1464 VDD VSS sg13g2_FILL8
XSTDFILL98_1472 VDD VSS sg13g2_FILL8
XSTDFILL98_1480 VDD VSS sg13g2_FILL8
XSTDFILL98_1488 VDD VSS sg13g2_FILL8
XSTDFILL98_1496 VDD VSS sg13g2_FILL8
XSTDFILL98_1504 VDD VSS sg13g2_FILL8
XSTDFILL98_1512 VDD VSS sg13g2_FILL8
XSTDFILL98_1520 VDD VSS sg13g2_FILL8
XSTDFILL98_1528 VDD VSS sg13g2_FILL2
XSTDFILL98_1530 VDD VSS sg13g2_FILL1
XSTDFILL99_0 VDD VSS sg13g2_FILL8
XSTDFILL99_8 VDD VSS sg13g2_FILL8
XSTDFILL99_16 VDD VSS sg13g2_FILL8
XSTDFILL99_24 VDD VSS sg13g2_FILL8
XSTDFILL99_32 VDD VSS sg13g2_FILL8
XSTDFILL99_40 VDD VSS sg13g2_FILL8
XSTDFILL99_48 VDD VSS sg13g2_FILL8
XSTDFILL99_56 VDD VSS sg13g2_FILL8
XSTDFILL99_64 VDD VSS sg13g2_FILL8
XSTDFILL99_72 VDD VSS sg13g2_FILL8
XSTDFILL99_80 VDD VSS sg13g2_FILL8
XSTDFILL99_88 VDD VSS sg13g2_FILL8
XSTDFILL99_96 VDD VSS sg13g2_FILL8
XSTDFILL99_104 VDD VSS sg13g2_FILL8
XSTDFILL99_112 VDD VSS sg13g2_FILL8
XSTDFILL99_120 VDD VSS sg13g2_FILL8
XSTDFILL99_128 VDD VSS sg13g2_FILL8
XSTDFILL99_136 VDD VSS sg13g2_FILL8
XSTDFILL99_144 VDD VSS sg13g2_FILL8
XSTDFILL99_152 VDD VSS sg13g2_FILL8
XSTDFILL99_160 VDD VSS sg13g2_FILL8
XSTDFILL99_168 VDD VSS sg13g2_FILL8
XSTDFILL99_176 VDD VSS sg13g2_FILL8
XSTDFILL99_184 VDD VSS sg13g2_FILL8
XSTDFILL99_192 VDD VSS sg13g2_FILL8
XSTDFILL99_200 VDD VSS sg13g2_FILL8
XSTDFILL99_208 VDD VSS sg13g2_FILL8
XSTDFILL99_216 VDD VSS sg13g2_FILL8
XSTDFILL99_224 VDD VSS sg13g2_FILL8
XSTDFILL99_232 VDD VSS sg13g2_FILL8
XSTDFILL99_240 VDD VSS sg13g2_FILL8
XSTDFILL99_248 VDD VSS sg13g2_FILL8
XSTDFILL99_256 VDD VSS sg13g2_FILL8
XSTDFILL99_264 VDD VSS sg13g2_FILL8
XSTDFILL99_272 VDD VSS sg13g2_FILL8
XSTDFILL99_280 VDD VSS sg13g2_FILL8
XSTDFILL99_288 VDD VSS sg13g2_FILL8
XSTDFILL99_296 VDD VSS sg13g2_FILL8
XSTDFILL99_304 VDD VSS sg13g2_FILL8
XSTDFILL99_312 VDD VSS sg13g2_FILL8
XSTDFILL99_320 VDD VSS sg13g2_FILL8
XSTDFILL99_328 VDD VSS sg13g2_FILL8
XSTDFILL99_336 VDD VSS sg13g2_FILL8
XSTDFILL99_344 VDD VSS sg13g2_FILL8
XSTDFILL99_352 VDD VSS sg13g2_FILL8
XSTDFILL99_360 VDD VSS sg13g2_FILL8
XSTDFILL99_368 VDD VSS sg13g2_FILL8
XSTDFILL99_376 VDD VSS sg13g2_FILL8
XSTDFILL99_384 VDD VSS sg13g2_FILL8
XSTDFILL99_392 VDD VSS sg13g2_FILL8
XSTDFILL99_400 VDD VSS sg13g2_FILL8
XSTDFILL99_408 VDD VSS sg13g2_FILL8
XSTDFILL99_416 VDD VSS sg13g2_FILL8
XSTDFILL99_424 VDD VSS sg13g2_FILL8
XSTDFILL99_432 VDD VSS sg13g2_FILL8
XSTDFILL99_440 VDD VSS sg13g2_FILL8
XSTDFILL99_448 VDD VSS sg13g2_FILL8
XSTDFILL99_456 VDD VSS sg13g2_FILL8
XSTDFILL99_464 VDD VSS sg13g2_FILL8
XSTDFILL99_472 VDD VSS sg13g2_FILL8
XSTDFILL99_480 VDD VSS sg13g2_FILL8
XSTDFILL99_488 VDD VSS sg13g2_FILL8
XSTDFILL99_496 VDD VSS sg13g2_FILL8
XSTDFILL99_504 VDD VSS sg13g2_FILL8
XSTDFILL99_512 VDD VSS sg13g2_FILL8
XSTDFILL99_520 VDD VSS sg13g2_FILL8
XSTDFILL99_528 VDD VSS sg13g2_FILL8
XSTDFILL99_536 VDD VSS sg13g2_FILL8
XSTDFILL99_544 VDD VSS sg13g2_FILL8
XSTDFILL99_552 VDD VSS sg13g2_FILL8
XSTDFILL99_560 VDD VSS sg13g2_FILL8
XSTDFILL99_568 VDD VSS sg13g2_FILL8
XSTDFILL99_576 VDD VSS sg13g2_FILL8
XSTDFILL99_584 VDD VSS sg13g2_FILL8
XSTDFILL99_592 VDD VSS sg13g2_FILL8
XSTDFILL99_600 VDD VSS sg13g2_FILL8
XSTDFILL99_608 VDD VSS sg13g2_FILL8
XSTDFILL99_616 VDD VSS sg13g2_FILL8
XSTDFILL99_624 VDD VSS sg13g2_FILL8
XSTDFILL99_632 VDD VSS sg13g2_FILL8
XSTDFILL99_640 VDD VSS sg13g2_FILL8
XSTDFILL99_648 VDD VSS sg13g2_FILL8
XSTDFILL99_656 VDD VSS sg13g2_FILL8
XSTDFILL99_664 VDD VSS sg13g2_FILL8
XSTDFILL99_672 VDD VSS sg13g2_FILL8
XSTDFILL99_680 VDD VSS sg13g2_FILL8
XSTDFILL99_688 VDD VSS sg13g2_FILL8
XSTDFILL99_696 VDD VSS sg13g2_FILL8
XSTDFILL99_704 VDD VSS sg13g2_FILL8
XSTDFILL99_712 VDD VSS sg13g2_FILL8
XSTDFILL99_720 VDD VSS sg13g2_FILL8
XSTDFILL99_728 VDD VSS sg13g2_FILL8
XSTDFILL99_736 VDD VSS sg13g2_FILL8
XSTDFILL99_744 VDD VSS sg13g2_FILL8
XSTDFILL99_752 VDD VSS sg13g2_FILL8
XSTDFILL99_760 VDD VSS sg13g2_FILL8
XSTDFILL99_768 VDD VSS sg13g2_FILL8
XSTDFILL99_776 VDD VSS sg13g2_FILL8
XSTDFILL99_784 VDD VSS sg13g2_FILL8
XSTDFILL99_792 VDD VSS sg13g2_FILL8
XSTDFILL99_800 VDD VSS sg13g2_FILL8
XSTDFILL99_808 VDD VSS sg13g2_FILL8
XSTDFILL99_816 VDD VSS sg13g2_FILL8
XSTDFILL99_824 VDD VSS sg13g2_FILL8
XSTDFILL99_832 VDD VSS sg13g2_FILL8
XSTDFILL99_840 VDD VSS sg13g2_FILL8
XSTDFILL99_848 VDD VSS sg13g2_FILL8
XSTDFILL99_856 VDD VSS sg13g2_FILL8
XSTDFILL99_864 VDD VSS sg13g2_FILL8
XSTDFILL99_872 VDD VSS sg13g2_FILL8
XSTDFILL99_880 VDD VSS sg13g2_FILL8
XSTDFILL99_888 VDD VSS sg13g2_FILL8
XSTDFILL99_896 VDD VSS sg13g2_FILL8
XSTDFILL99_904 VDD VSS sg13g2_FILL8
XSTDFILL99_912 VDD VSS sg13g2_FILL8
XSTDFILL99_920 VDD VSS sg13g2_FILL8
XSTDFILL99_928 VDD VSS sg13g2_FILL8
XSTDFILL99_936 VDD VSS sg13g2_FILL8
XSTDFILL99_944 VDD VSS sg13g2_FILL8
XSTDFILL99_952 VDD VSS sg13g2_FILL8
XSTDFILL99_960 VDD VSS sg13g2_FILL8
XSTDFILL99_968 VDD VSS sg13g2_FILL8
XSTDFILL99_976 VDD VSS sg13g2_FILL8
XSTDFILL99_984 VDD VSS sg13g2_FILL8
XSTDFILL99_992 VDD VSS sg13g2_FILL8
XSTDFILL99_1000 VDD VSS sg13g2_FILL8
XSTDFILL99_1008 VDD VSS sg13g2_FILL8
XSTDFILL99_1016 VDD VSS sg13g2_FILL8
XSTDFILL99_1024 VDD VSS sg13g2_FILL8
XSTDFILL99_1032 VDD VSS sg13g2_FILL8
XSTDFILL99_1040 VDD VSS sg13g2_FILL8
XSTDFILL99_1048 VDD VSS sg13g2_FILL8
XSTDFILL99_1056 VDD VSS sg13g2_FILL8
XSTDFILL99_1064 VDD VSS sg13g2_FILL8
XSTDFILL99_1072 VDD VSS sg13g2_FILL8
XSTDFILL99_1080 VDD VSS sg13g2_FILL8
XSTDFILL99_1088 VDD VSS sg13g2_FILL8
XSTDFILL99_1096 VDD VSS sg13g2_FILL8
XSTDFILL99_1104 VDD VSS sg13g2_FILL8
XSTDFILL99_1112 VDD VSS sg13g2_FILL8
XSTDFILL99_1120 VDD VSS sg13g2_FILL8
XSTDFILL99_1128 VDD VSS sg13g2_FILL8
XSTDFILL99_1136 VDD VSS sg13g2_FILL8
XSTDFILL99_1144 VDD VSS sg13g2_FILL8
XSTDFILL99_1152 VDD VSS sg13g2_FILL8
XSTDFILL99_1160 VDD VSS sg13g2_FILL8
XSTDFILL99_1168 VDD VSS sg13g2_FILL8
XSTDFILL99_1176 VDD VSS sg13g2_FILL8
XSTDFILL99_1184 VDD VSS sg13g2_FILL8
XSTDFILL99_1192 VDD VSS sg13g2_FILL8
XSTDFILL99_1200 VDD VSS sg13g2_FILL8
XSTDFILL99_1208 VDD VSS sg13g2_FILL8
XSTDFILL99_1216 VDD VSS sg13g2_FILL8
XSTDFILL99_1224 VDD VSS sg13g2_FILL8
XSTDFILL99_1232 VDD VSS sg13g2_FILL8
XSTDFILL99_1240 VDD VSS sg13g2_FILL8
XSTDFILL99_1248 VDD VSS sg13g2_FILL8
XSTDFILL99_1256 VDD VSS sg13g2_FILL8
XSTDFILL99_1264 VDD VSS sg13g2_FILL8
XSTDFILL99_1272 VDD VSS sg13g2_FILL8
XSTDFILL99_1280 VDD VSS sg13g2_FILL8
XSTDFILL99_1288 VDD VSS sg13g2_FILL8
XSTDFILL99_1296 VDD VSS sg13g2_FILL8
XSTDFILL99_1304 VDD VSS sg13g2_FILL8
XSTDFILL99_1312 VDD VSS sg13g2_FILL8
XSTDFILL99_1320 VDD VSS sg13g2_FILL8
XSTDFILL99_1328 VDD VSS sg13g2_FILL8
XSTDFILL99_1336 VDD VSS sg13g2_FILL8
XSTDFILL99_1344 VDD VSS sg13g2_FILL8
XSTDFILL99_1352 VDD VSS sg13g2_FILL8
XSTDFILL99_1360 VDD VSS sg13g2_FILL8
XSTDFILL99_1368 VDD VSS sg13g2_FILL8
XSTDFILL99_1376 VDD VSS sg13g2_FILL8
XSTDFILL99_1384 VDD VSS sg13g2_FILL8
XSTDFILL99_1392 VDD VSS sg13g2_FILL8
XSTDFILL99_1400 VDD VSS sg13g2_FILL8
XSTDFILL99_1408 VDD VSS sg13g2_FILL8
XSTDFILL99_1416 VDD VSS sg13g2_FILL8
XSTDFILL99_1424 VDD VSS sg13g2_FILL8
XSTDFILL99_1432 VDD VSS sg13g2_FILL8
XSTDFILL99_1440 VDD VSS sg13g2_FILL8
XSTDFILL99_1448 VDD VSS sg13g2_FILL8
XSTDFILL99_1456 VDD VSS sg13g2_FILL8
XSTDFILL99_1464 VDD VSS sg13g2_FILL8
XSTDFILL99_1472 VDD VSS sg13g2_FILL8
XSTDFILL99_1480 VDD VSS sg13g2_FILL8
XSTDFILL99_1488 VDD VSS sg13g2_FILL8
XSTDFILL99_1496 VDD VSS sg13g2_FILL8
XSTDFILL99_1504 VDD VSS sg13g2_FILL8
XSTDFILL99_1512 VDD VSS sg13g2_FILL8
XSTDFILL99_1520 VDD VSS sg13g2_FILL8
XSTDFILL99_1528 VDD VSS sg13g2_FILL2
XSTDFILL99_1530 VDD VSS sg13g2_FILL1
XSTDFILL100_0 VDD VSS sg13g2_FILL8
XSTDFILL100_8 VDD VSS sg13g2_FILL8
XSTDFILL100_16 VDD VSS sg13g2_FILL8
XSTDFILL100_24 VDD VSS sg13g2_FILL8
XSTDFILL100_32 VDD VSS sg13g2_FILL8
XSTDFILL100_40 VDD VSS sg13g2_FILL8
XSTDFILL100_48 VDD VSS sg13g2_FILL8
XSTDFILL100_56 VDD VSS sg13g2_FILL8
XSTDFILL100_64 VDD VSS sg13g2_FILL8
XSTDFILL100_72 VDD VSS sg13g2_FILL8
XSTDFILL100_80 VDD VSS sg13g2_FILL8
XSTDFILL100_88 VDD VSS sg13g2_FILL8
XSTDFILL100_96 VDD VSS sg13g2_FILL8
XSTDFILL100_104 VDD VSS sg13g2_FILL8
XSTDFILL100_112 VDD VSS sg13g2_FILL8
XSTDFILL100_120 VDD VSS sg13g2_FILL8
XSTDFILL100_128 VDD VSS sg13g2_FILL8
XSTDFILL100_136 VDD VSS sg13g2_FILL8
XSTDFILL100_144 VDD VSS sg13g2_FILL8
XSTDFILL100_152 VDD VSS sg13g2_FILL8
XSTDFILL100_160 VDD VSS sg13g2_FILL8
XSTDFILL100_168 VDD VSS sg13g2_FILL8
XSTDFILL100_176 VDD VSS sg13g2_FILL8
XSTDFILL100_184 VDD VSS sg13g2_FILL8
XSTDFILL100_192 VDD VSS sg13g2_FILL8
XSTDFILL100_200 VDD VSS sg13g2_FILL8
XSTDFILL100_208 VDD VSS sg13g2_FILL8
XSTDFILL100_216 VDD VSS sg13g2_FILL8
XSTDFILL100_224 VDD VSS sg13g2_FILL8
XSTDFILL100_232 VDD VSS sg13g2_FILL8
XSTDFILL100_240 VDD VSS sg13g2_FILL8
XSTDFILL100_248 VDD VSS sg13g2_FILL8
XSTDFILL100_256 VDD VSS sg13g2_FILL8
XSTDFILL100_264 VDD VSS sg13g2_FILL8
XSTDFILL100_272 VDD VSS sg13g2_FILL8
XSTDFILL100_280 VDD VSS sg13g2_FILL8
XSTDFILL100_288 VDD VSS sg13g2_FILL8
XSTDFILL100_296 VDD VSS sg13g2_FILL8
XSTDFILL100_304 VDD VSS sg13g2_FILL8
XSTDFILL100_312 VDD VSS sg13g2_FILL8
XSTDFILL100_320 VDD VSS sg13g2_FILL8
XSTDFILL100_328 VDD VSS sg13g2_FILL8
XSTDFILL100_336 VDD VSS sg13g2_FILL8
XSTDFILL100_344 VDD VSS sg13g2_FILL8
XSTDFILL100_352 VDD VSS sg13g2_FILL8
XSTDFILL100_360 VDD VSS sg13g2_FILL8
XSTDFILL100_368 VDD VSS sg13g2_FILL8
XSTDFILL100_376 VDD VSS sg13g2_FILL8
XSTDFILL100_384 VDD VSS sg13g2_FILL8
XSTDFILL100_392 VDD VSS sg13g2_FILL8
XSTDFILL100_400 VDD VSS sg13g2_FILL8
XSTDFILL100_408 VDD VSS sg13g2_FILL8
XSTDFILL100_416 VDD VSS sg13g2_FILL8
XSTDFILL100_424 VDD VSS sg13g2_FILL8
XSTDFILL100_432 VDD VSS sg13g2_FILL8
XSTDFILL100_440 VDD VSS sg13g2_FILL8
XSTDFILL100_448 VDD VSS sg13g2_FILL8
XSTDFILL100_456 VDD VSS sg13g2_FILL8
XSTDFILL100_464 VDD VSS sg13g2_FILL8
XSTDFILL100_472 VDD VSS sg13g2_FILL8
XSTDFILL100_480 VDD VSS sg13g2_FILL8
XSTDFILL100_488 VDD VSS sg13g2_FILL8
XSTDFILL100_496 VDD VSS sg13g2_FILL8
XSTDFILL100_504 VDD VSS sg13g2_FILL8
XSTDFILL100_512 VDD VSS sg13g2_FILL8
XSTDFILL100_520 VDD VSS sg13g2_FILL8
XSTDFILL100_528 VDD VSS sg13g2_FILL8
XSTDFILL100_536 VDD VSS sg13g2_FILL8
XSTDFILL100_544 VDD VSS sg13g2_FILL8
XSTDFILL100_552 VDD VSS sg13g2_FILL8
XSTDFILL100_560 VDD VSS sg13g2_FILL8
XSTDFILL100_568 VDD VSS sg13g2_FILL8
XSTDFILL100_576 VDD VSS sg13g2_FILL8
XSTDFILL100_584 VDD VSS sg13g2_FILL8
XSTDFILL100_592 VDD VSS sg13g2_FILL8
XSTDFILL100_600 VDD VSS sg13g2_FILL8
XSTDFILL100_608 VDD VSS sg13g2_FILL8
XSTDFILL100_616 VDD VSS sg13g2_FILL8
XSTDFILL100_624 VDD VSS sg13g2_FILL8
XSTDFILL100_632 VDD VSS sg13g2_FILL8
XSTDFILL100_640 VDD VSS sg13g2_FILL8
XSTDFILL100_648 VDD VSS sg13g2_FILL8
XSTDFILL100_656 VDD VSS sg13g2_FILL8
XSTDFILL100_664 VDD VSS sg13g2_FILL8
XSTDFILL100_672 VDD VSS sg13g2_FILL8
XSTDFILL100_680 VDD VSS sg13g2_FILL8
XSTDFILL100_688 VDD VSS sg13g2_FILL8
XSTDFILL100_696 VDD VSS sg13g2_FILL8
XSTDFILL100_704 VDD VSS sg13g2_FILL8
XSTDFILL100_712 VDD VSS sg13g2_FILL8
XSTDFILL100_720 VDD VSS sg13g2_FILL8
XSTDFILL100_728 VDD VSS sg13g2_FILL8
XSTDFILL100_736 VDD VSS sg13g2_FILL8
XSTDFILL100_744 VDD VSS sg13g2_FILL8
XSTDFILL100_752 VDD VSS sg13g2_FILL8
XSTDFILL100_760 VDD VSS sg13g2_FILL8
XSTDFILL100_768 VDD VSS sg13g2_FILL8
XSTDFILL100_776 VDD VSS sg13g2_FILL8
XSTDFILL100_784 VDD VSS sg13g2_FILL8
XSTDFILL100_792 VDD VSS sg13g2_FILL8
XSTDFILL100_800 VDD VSS sg13g2_FILL8
XSTDFILL100_808 VDD VSS sg13g2_FILL8
XSTDFILL100_816 VDD VSS sg13g2_FILL8
XSTDFILL100_824 VDD VSS sg13g2_FILL8
XSTDFILL100_832 VDD VSS sg13g2_FILL8
XSTDFILL100_840 VDD VSS sg13g2_FILL8
XSTDFILL100_848 VDD VSS sg13g2_FILL8
XSTDFILL100_856 VDD VSS sg13g2_FILL8
XSTDFILL100_864 VDD VSS sg13g2_FILL8
XSTDFILL100_872 VDD VSS sg13g2_FILL8
XSTDFILL100_880 VDD VSS sg13g2_FILL8
XSTDFILL100_888 VDD VSS sg13g2_FILL8
XSTDFILL100_896 VDD VSS sg13g2_FILL8
XSTDFILL100_904 VDD VSS sg13g2_FILL8
XSTDFILL100_912 VDD VSS sg13g2_FILL8
XSTDFILL100_920 VDD VSS sg13g2_FILL8
XSTDFILL100_928 VDD VSS sg13g2_FILL8
XSTDFILL100_936 VDD VSS sg13g2_FILL8
XSTDFILL100_944 VDD VSS sg13g2_FILL8
XSTDFILL100_952 VDD VSS sg13g2_FILL8
XSTDFILL100_960 VDD VSS sg13g2_FILL8
XSTDFILL100_968 VDD VSS sg13g2_FILL8
XSTDFILL100_976 VDD VSS sg13g2_FILL8
XSTDFILL100_984 VDD VSS sg13g2_FILL8
XSTDFILL100_992 VDD VSS sg13g2_FILL8
XSTDFILL100_1000 VDD VSS sg13g2_FILL8
XSTDFILL100_1008 VDD VSS sg13g2_FILL8
XSTDFILL100_1016 VDD VSS sg13g2_FILL8
XSTDFILL100_1024 VDD VSS sg13g2_FILL8
XSTDFILL100_1032 VDD VSS sg13g2_FILL8
XSTDFILL100_1040 VDD VSS sg13g2_FILL8
XSTDFILL100_1048 VDD VSS sg13g2_FILL8
XSTDFILL100_1056 VDD VSS sg13g2_FILL8
XSTDFILL100_1064 VDD VSS sg13g2_FILL8
XSTDFILL100_1072 VDD VSS sg13g2_FILL8
XSTDFILL100_1080 VDD VSS sg13g2_FILL8
XSTDFILL100_1088 VDD VSS sg13g2_FILL8
XSTDFILL100_1096 VDD VSS sg13g2_FILL8
XSTDFILL100_1104 VDD VSS sg13g2_FILL8
XSTDFILL100_1112 VDD VSS sg13g2_FILL8
XSTDFILL100_1120 VDD VSS sg13g2_FILL8
XSTDFILL100_1128 VDD VSS sg13g2_FILL8
XSTDFILL100_1136 VDD VSS sg13g2_FILL8
XSTDFILL100_1144 VDD VSS sg13g2_FILL8
XSTDFILL100_1152 VDD VSS sg13g2_FILL8
XSTDFILL100_1160 VDD VSS sg13g2_FILL8
XSTDFILL100_1168 VDD VSS sg13g2_FILL8
XSTDFILL100_1176 VDD VSS sg13g2_FILL8
XSTDFILL100_1184 VDD VSS sg13g2_FILL8
XSTDFILL100_1192 VDD VSS sg13g2_FILL8
XSTDFILL100_1200 VDD VSS sg13g2_FILL8
XSTDFILL100_1208 VDD VSS sg13g2_FILL8
XSTDFILL100_1216 VDD VSS sg13g2_FILL8
XSTDFILL100_1224 VDD VSS sg13g2_FILL8
XSTDFILL100_1232 VDD VSS sg13g2_FILL8
XSTDFILL100_1240 VDD VSS sg13g2_FILL8
XSTDFILL100_1248 VDD VSS sg13g2_FILL8
XSTDFILL100_1256 VDD VSS sg13g2_FILL8
XSTDFILL100_1264 VDD VSS sg13g2_FILL8
XSTDFILL100_1272 VDD VSS sg13g2_FILL8
XSTDFILL100_1280 VDD VSS sg13g2_FILL8
XSTDFILL100_1288 VDD VSS sg13g2_FILL8
XSTDFILL100_1296 VDD VSS sg13g2_FILL8
XSTDFILL100_1304 VDD VSS sg13g2_FILL8
XSTDFILL100_1312 VDD VSS sg13g2_FILL8
XSTDFILL100_1320 VDD VSS sg13g2_FILL8
XSTDFILL100_1328 VDD VSS sg13g2_FILL8
XSTDFILL100_1336 VDD VSS sg13g2_FILL8
XSTDFILL100_1344 VDD VSS sg13g2_FILL8
XSTDFILL100_1352 VDD VSS sg13g2_FILL8
XSTDFILL100_1360 VDD VSS sg13g2_FILL8
XSTDFILL100_1368 VDD VSS sg13g2_FILL8
XSTDFILL100_1376 VDD VSS sg13g2_FILL8
XSTDFILL100_1384 VDD VSS sg13g2_FILL8
XSTDFILL100_1392 VDD VSS sg13g2_FILL8
XSTDFILL100_1400 VDD VSS sg13g2_FILL8
XSTDFILL100_1408 VDD VSS sg13g2_FILL8
XSTDFILL100_1416 VDD VSS sg13g2_FILL8
XSTDFILL100_1424 VDD VSS sg13g2_FILL8
XSTDFILL100_1432 VDD VSS sg13g2_FILL8
XSTDFILL100_1440 VDD VSS sg13g2_FILL8
XSTDFILL100_1448 VDD VSS sg13g2_FILL8
XSTDFILL100_1456 VDD VSS sg13g2_FILL8
XSTDFILL100_1464 VDD VSS sg13g2_FILL8
XSTDFILL100_1472 VDD VSS sg13g2_FILL8
XSTDFILL100_1480 VDD VSS sg13g2_FILL8
XSTDFILL100_1488 VDD VSS sg13g2_FILL8
XSTDFILL100_1496 VDD VSS sg13g2_FILL8
XSTDFILL100_1504 VDD VSS sg13g2_FILL8
XSTDFILL100_1512 VDD VSS sg13g2_FILL8
XSTDFILL100_1520 VDD VSS sg13g2_FILL8
XSTDFILL100_1528 VDD VSS sg13g2_FILL2
XSTDFILL100_1530 VDD VSS sg13g2_FILL1
XSTDFILL101_0 VDD VSS sg13g2_FILL8
XSTDFILL101_8 VDD VSS sg13g2_FILL8
XSTDFILL101_16 VDD VSS sg13g2_FILL8
XSTDFILL101_24 VDD VSS sg13g2_FILL8
XSTDFILL101_32 VDD VSS sg13g2_FILL8
XSTDFILL101_40 VDD VSS sg13g2_FILL8
XSTDFILL101_48 VDD VSS sg13g2_FILL8
XSTDFILL101_56 VDD VSS sg13g2_FILL8
XSTDFILL101_64 VDD VSS sg13g2_FILL8
XSTDFILL101_72 VDD VSS sg13g2_FILL8
XSTDFILL101_80 VDD VSS sg13g2_FILL8
XSTDFILL101_88 VDD VSS sg13g2_FILL8
XSTDFILL101_96 VDD VSS sg13g2_FILL8
XSTDFILL101_104 VDD VSS sg13g2_FILL8
XSTDFILL101_112 VDD VSS sg13g2_FILL8
XSTDFILL101_120 VDD VSS sg13g2_FILL8
XSTDFILL101_128 VDD VSS sg13g2_FILL8
XSTDFILL101_136 VDD VSS sg13g2_FILL8
XSTDFILL101_144 VDD VSS sg13g2_FILL8
XSTDFILL101_152 VDD VSS sg13g2_FILL8
XSTDFILL101_160 VDD VSS sg13g2_FILL8
XSTDFILL101_168 VDD VSS sg13g2_FILL8
XSTDFILL101_176 VDD VSS sg13g2_FILL8
XSTDFILL101_184 VDD VSS sg13g2_FILL8
XSTDFILL101_192 VDD VSS sg13g2_FILL8
XSTDFILL101_200 VDD VSS sg13g2_FILL8
XSTDFILL101_208 VDD VSS sg13g2_FILL8
XSTDFILL101_216 VDD VSS sg13g2_FILL8
XSTDFILL101_224 VDD VSS sg13g2_FILL8
XSTDFILL101_232 VDD VSS sg13g2_FILL8
XSTDFILL101_240 VDD VSS sg13g2_FILL8
XSTDFILL101_248 VDD VSS sg13g2_FILL8
XSTDFILL101_256 VDD VSS sg13g2_FILL8
XSTDFILL101_264 VDD VSS sg13g2_FILL8
XSTDFILL101_272 VDD VSS sg13g2_FILL8
XSTDFILL101_280 VDD VSS sg13g2_FILL8
XSTDFILL101_288 VDD VSS sg13g2_FILL8
XSTDFILL101_296 VDD VSS sg13g2_FILL8
XSTDFILL101_304 VDD VSS sg13g2_FILL8
XSTDFILL101_312 VDD VSS sg13g2_FILL8
XSTDFILL101_320 VDD VSS sg13g2_FILL8
XSTDFILL101_328 VDD VSS sg13g2_FILL8
XSTDFILL101_336 VDD VSS sg13g2_FILL8
XSTDFILL101_344 VDD VSS sg13g2_FILL8
XSTDFILL101_352 VDD VSS sg13g2_FILL8
XSTDFILL101_360 VDD VSS sg13g2_FILL8
XSTDFILL101_368 VDD VSS sg13g2_FILL8
XSTDFILL101_376 VDD VSS sg13g2_FILL8
XSTDFILL101_384 VDD VSS sg13g2_FILL8
XSTDFILL101_392 VDD VSS sg13g2_FILL8
XSTDFILL101_400 VDD VSS sg13g2_FILL8
XSTDFILL101_408 VDD VSS sg13g2_FILL8
XSTDFILL101_416 VDD VSS sg13g2_FILL8
XSTDFILL101_424 VDD VSS sg13g2_FILL8
XSTDFILL101_432 VDD VSS sg13g2_FILL8
XSTDFILL101_440 VDD VSS sg13g2_FILL8
XSTDFILL101_448 VDD VSS sg13g2_FILL8
XSTDFILL101_456 VDD VSS sg13g2_FILL8
XSTDFILL101_464 VDD VSS sg13g2_FILL8
XSTDFILL101_472 VDD VSS sg13g2_FILL8
XSTDFILL101_480 VDD VSS sg13g2_FILL8
XSTDFILL101_488 VDD VSS sg13g2_FILL8
XSTDFILL101_496 VDD VSS sg13g2_FILL8
XSTDFILL101_504 VDD VSS sg13g2_FILL8
XSTDFILL101_512 VDD VSS sg13g2_FILL8
XSTDFILL101_520 VDD VSS sg13g2_FILL8
XSTDFILL101_528 VDD VSS sg13g2_FILL8
XSTDFILL101_536 VDD VSS sg13g2_FILL8
XSTDFILL101_544 VDD VSS sg13g2_FILL8
XSTDFILL101_552 VDD VSS sg13g2_FILL8
XSTDFILL101_560 VDD VSS sg13g2_FILL8
XSTDFILL101_568 VDD VSS sg13g2_FILL8
XSTDFILL101_576 VDD VSS sg13g2_FILL8
XSTDFILL101_584 VDD VSS sg13g2_FILL8
XSTDFILL101_592 VDD VSS sg13g2_FILL8
XSTDFILL101_600 VDD VSS sg13g2_FILL8
XSTDFILL101_608 VDD VSS sg13g2_FILL8
XSTDFILL101_616 VDD VSS sg13g2_FILL8
XSTDFILL101_624 VDD VSS sg13g2_FILL8
XSTDFILL101_632 VDD VSS sg13g2_FILL8
XSTDFILL101_640 VDD VSS sg13g2_FILL8
XSTDFILL101_648 VDD VSS sg13g2_FILL8
XSTDFILL101_656 VDD VSS sg13g2_FILL8
XSTDFILL101_664 VDD VSS sg13g2_FILL8
XSTDFILL101_672 VDD VSS sg13g2_FILL8
XSTDFILL101_680 VDD VSS sg13g2_FILL8
XSTDFILL101_688 VDD VSS sg13g2_FILL8
XSTDFILL101_696 VDD VSS sg13g2_FILL8
XSTDFILL101_704 VDD VSS sg13g2_FILL8
XSTDFILL101_712 VDD VSS sg13g2_FILL8
XSTDFILL101_720 VDD VSS sg13g2_FILL8
XSTDFILL101_728 VDD VSS sg13g2_FILL8
XSTDFILL101_736 VDD VSS sg13g2_FILL8
XSTDFILL101_744 VDD VSS sg13g2_FILL8
XSTDFILL101_752 VDD VSS sg13g2_FILL8
XSTDFILL101_760 VDD VSS sg13g2_FILL8
XSTDFILL101_768 VDD VSS sg13g2_FILL8
XSTDFILL101_776 VDD VSS sg13g2_FILL8
XSTDFILL101_784 VDD VSS sg13g2_FILL8
XSTDFILL101_792 VDD VSS sg13g2_FILL8
XSTDFILL101_800 VDD VSS sg13g2_FILL8
XSTDFILL101_808 VDD VSS sg13g2_FILL8
XSTDFILL101_816 VDD VSS sg13g2_FILL8
XSTDFILL101_824 VDD VSS sg13g2_FILL8
XSTDFILL101_832 VDD VSS sg13g2_FILL8
XSTDFILL101_840 VDD VSS sg13g2_FILL8
XSTDFILL101_848 VDD VSS sg13g2_FILL8
XSTDFILL101_856 VDD VSS sg13g2_FILL8
XSTDFILL101_864 VDD VSS sg13g2_FILL8
XSTDFILL101_872 VDD VSS sg13g2_FILL8
XSTDFILL101_880 VDD VSS sg13g2_FILL8
XSTDFILL101_888 VDD VSS sg13g2_FILL8
XSTDFILL101_896 VDD VSS sg13g2_FILL8
XSTDFILL101_904 VDD VSS sg13g2_FILL8
XSTDFILL101_912 VDD VSS sg13g2_FILL8
XSTDFILL101_920 VDD VSS sg13g2_FILL8
XSTDFILL101_928 VDD VSS sg13g2_FILL8
XSTDFILL101_936 VDD VSS sg13g2_FILL8
XSTDFILL101_944 VDD VSS sg13g2_FILL8
XSTDFILL101_952 VDD VSS sg13g2_FILL8
XSTDFILL101_960 VDD VSS sg13g2_FILL8
XSTDFILL101_968 VDD VSS sg13g2_FILL8
XSTDFILL101_976 VDD VSS sg13g2_FILL8
XSTDFILL101_984 VDD VSS sg13g2_FILL8
XSTDFILL101_992 VDD VSS sg13g2_FILL8
XSTDFILL101_1000 VDD VSS sg13g2_FILL8
XSTDFILL101_1008 VDD VSS sg13g2_FILL8
XSTDFILL101_1016 VDD VSS sg13g2_FILL8
XSTDFILL101_1024 VDD VSS sg13g2_FILL8
XSTDFILL101_1032 VDD VSS sg13g2_FILL8
XSTDFILL101_1040 VDD VSS sg13g2_FILL8
XSTDFILL101_1048 VDD VSS sg13g2_FILL8
XSTDFILL101_1056 VDD VSS sg13g2_FILL8
XSTDFILL101_1064 VDD VSS sg13g2_FILL8
XSTDFILL101_1072 VDD VSS sg13g2_FILL8
XSTDFILL101_1080 VDD VSS sg13g2_FILL8
XSTDFILL101_1088 VDD VSS sg13g2_FILL8
XSTDFILL101_1096 VDD VSS sg13g2_FILL8
XSTDFILL101_1104 VDD VSS sg13g2_FILL8
XSTDFILL101_1112 VDD VSS sg13g2_FILL8
XSTDFILL101_1120 VDD VSS sg13g2_FILL8
XSTDFILL101_1128 VDD VSS sg13g2_FILL8
XSTDFILL101_1136 VDD VSS sg13g2_FILL8
XSTDFILL101_1144 VDD VSS sg13g2_FILL8
XSTDFILL101_1152 VDD VSS sg13g2_FILL8
XSTDFILL101_1160 VDD VSS sg13g2_FILL8
XSTDFILL101_1168 VDD VSS sg13g2_FILL8
XSTDFILL101_1176 VDD VSS sg13g2_FILL8
XSTDFILL101_1184 VDD VSS sg13g2_FILL8
XSTDFILL101_1192 VDD VSS sg13g2_FILL8
XSTDFILL101_1200 VDD VSS sg13g2_FILL8
XSTDFILL101_1208 VDD VSS sg13g2_FILL8
XSTDFILL101_1216 VDD VSS sg13g2_FILL8
XSTDFILL101_1224 VDD VSS sg13g2_FILL8
XSTDFILL101_1232 VDD VSS sg13g2_FILL8
XSTDFILL101_1240 VDD VSS sg13g2_FILL8
XSTDFILL101_1248 VDD VSS sg13g2_FILL8
XSTDFILL101_1256 VDD VSS sg13g2_FILL8
XSTDFILL101_1264 VDD VSS sg13g2_FILL8
XSTDFILL101_1272 VDD VSS sg13g2_FILL8
XSTDFILL101_1280 VDD VSS sg13g2_FILL8
XSTDFILL101_1288 VDD VSS sg13g2_FILL8
XSTDFILL101_1296 VDD VSS sg13g2_FILL8
XSTDFILL101_1304 VDD VSS sg13g2_FILL8
XSTDFILL101_1312 VDD VSS sg13g2_FILL8
XSTDFILL101_1320 VDD VSS sg13g2_FILL8
XSTDFILL101_1328 VDD VSS sg13g2_FILL8
XSTDFILL101_1336 VDD VSS sg13g2_FILL8
XSTDFILL101_1344 VDD VSS sg13g2_FILL8
XSTDFILL101_1352 VDD VSS sg13g2_FILL8
XSTDFILL101_1360 VDD VSS sg13g2_FILL8
XSTDFILL101_1368 VDD VSS sg13g2_FILL8
XSTDFILL101_1376 VDD VSS sg13g2_FILL8
XSTDFILL101_1384 VDD VSS sg13g2_FILL8
XSTDFILL101_1392 VDD VSS sg13g2_FILL8
XSTDFILL101_1400 VDD VSS sg13g2_FILL8
XSTDFILL101_1408 VDD VSS sg13g2_FILL8
XSTDFILL101_1416 VDD VSS sg13g2_FILL8
XSTDFILL101_1424 VDD VSS sg13g2_FILL8
XSTDFILL101_1432 VDD VSS sg13g2_FILL8
XSTDFILL101_1440 VDD VSS sg13g2_FILL8
XSTDFILL101_1448 VDD VSS sg13g2_FILL8
XSTDFILL101_1456 VDD VSS sg13g2_FILL8
XSTDFILL101_1464 VDD VSS sg13g2_FILL8
XSTDFILL101_1472 VDD VSS sg13g2_FILL8
XSTDFILL101_1480 VDD VSS sg13g2_FILL8
XSTDFILL101_1488 VDD VSS sg13g2_FILL8
XSTDFILL101_1496 VDD VSS sg13g2_FILL8
XSTDFILL101_1504 VDD VSS sg13g2_FILL8
XSTDFILL101_1512 VDD VSS sg13g2_FILL8
XSTDFILL101_1520 VDD VSS sg13g2_FILL8
XSTDFILL101_1528 VDD VSS sg13g2_FILL2
XSTDFILL101_1530 VDD VSS sg13g2_FILL1
XSTDFILL102_0 VDD VSS sg13g2_FILL8
XSTDFILL102_8 VDD VSS sg13g2_FILL8
XSTDFILL102_16 VDD VSS sg13g2_FILL8
XSTDFILL102_24 VDD VSS sg13g2_FILL8
XSTDFILL102_32 VDD VSS sg13g2_FILL8
XSTDFILL102_40 VDD VSS sg13g2_FILL8
XSTDFILL102_48 VDD VSS sg13g2_FILL8
XSTDFILL102_56 VDD VSS sg13g2_FILL8
XSTDFILL102_64 VDD VSS sg13g2_FILL8
XSTDFILL102_72 VDD VSS sg13g2_FILL8
XSTDFILL102_80 VDD VSS sg13g2_FILL8
XSTDFILL102_88 VDD VSS sg13g2_FILL8
XSTDFILL102_96 VDD VSS sg13g2_FILL8
XSTDFILL102_104 VDD VSS sg13g2_FILL8
XSTDFILL102_112 VDD VSS sg13g2_FILL8
XSTDFILL102_120 VDD VSS sg13g2_FILL8
XSTDFILL102_128 VDD VSS sg13g2_FILL8
XSTDFILL102_136 VDD VSS sg13g2_FILL8
XSTDFILL102_144 VDD VSS sg13g2_FILL8
XSTDFILL102_152 VDD VSS sg13g2_FILL8
XSTDFILL102_160 VDD VSS sg13g2_FILL8
XSTDFILL102_168 VDD VSS sg13g2_FILL8
XSTDFILL102_176 VDD VSS sg13g2_FILL8
XSTDFILL102_184 VDD VSS sg13g2_FILL8
XSTDFILL102_192 VDD VSS sg13g2_FILL8
XSTDFILL102_200 VDD VSS sg13g2_FILL8
XSTDFILL102_208 VDD VSS sg13g2_FILL8
XSTDFILL102_216 VDD VSS sg13g2_FILL8
XSTDFILL102_224 VDD VSS sg13g2_FILL8
XSTDFILL102_232 VDD VSS sg13g2_FILL8
XSTDFILL102_240 VDD VSS sg13g2_FILL8
XSTDFILL102_248 VDD VSS sg13g2_FILL8
XSTDFILL102_256 VDD VSS sg13g2_FILL8
XSTDFILL102_264 VDD VSS sg13g2_FILL8
XSTDFILL102_272 VDD VSS sg13g2_FILL8
XSTDFILL102_280 VDD VSS sg13g2_FILL8
XSTDFILL102_288 VDD VSS sg13g2_FILL8
XSTDFILL102_296 VDD VSS sg13g2_FILL8
XSTDFILL102_304 VDD VSS sg13g2_FILL8
XSTDFILL102_312 VDD VSS sg13g2_FILL8
XSTDFILL102_320 VDD VSS sg13g2_FILL8
XSTDFILL102_328 VDD VSS sg13g2_FILL8
XSTDFILL102_336 VDD VSS sg13g2_FILL8
XSTDFILL102_344 VDD VSS sg13g2_FILL8
XSTDFILL102_352 VDD VSS sg13g2_FILL8
XSTDFILL102_360 VDD VSS sg13g2_FILL8
XSTDFILL102_368 VDD VSS sg13g2_FILL8
XSTDFILL102_376 VDD VSS sg13g2_FILL8
XSTDFILL102_384 VDD VSS sg13g2_FILL8
XSTDFILL102_392 VDD VSS sg13g2_FILL8
XSTDFILL102_400 VDD VSS sg13g2_FILL8
XSTDFILL102_408 VDD VSS sg13g2_FILL8
XSTDFILL102_416 VDD VSS sg13g2_FILL8
XSTDFILL102_424 VDD VSS sg13g2_FILL8
XSTDFILL102_432 VDD VSS sg13g2_FILL8
XSTDFILL102_440 VDD VSS sg13g2_FILL8
XSTDFILL102_448 VDD VSS sg13g2_FILL8
XSTDFILL102_456 VDD VSS sg13g2_FILL8
XSTDFILL102_464 VDD VSS sg13g2_FILL8
XSTDFILL102_472 VDD VSS sg13g2_FILL8
XSTDFILL102_480 VDD VSS sg13g2_FILL8
XSTDFILL102_488 VDD VSS sg13g2_FILL8
XSTDFILL102_496 VDD VSS sg13g2_FILL8
XSTDFILL102_504 VDD VSS sg13g2_FILL8
XSTDFILL102_512 VDD VSS sg13g2_FILL8
XSTDFILL102_520 VDD VSS sg13g2_FILL8
XSTDFILL102_528 VDD VSS sg13g2_FILL8
XSTDFILL102_536 VDD VSS sg13g2_FILL8
XSTDFILL102_544 VDD VSS sg13g2_FILL8
XSTDFILL102_552 VDD VSS sg13g2_FILL8
XSTDFILL102_560 VDD VSS sg13g2_FILL8
XSTDFILL102_568 VDD VSS sg13g2_FILL8
XSTDFILL102_576 VDD VSS sg13g2_FILL8
XSTDFILL102_584 VDD VSS sg13g2_FILL8
XSTDFILL102_592 VDD VSS sg13g2_FILL8
XSTDFILL102_600 VDD VSS sg13g2_FILL8
XSTDFILL102_608 VDD VSS sg13g2_FILL8
XSTDFILL102_616 VDD VSS sg13g2_FILL8
XSTDFILL102_624 VDD VSS sg13g2_FILL8
XSTDFILL102_632 VDD VSS sg13g2_FILL8
XSTDFILL102_640 VDD VSS sg13g2_FILL8
XSTDFILL102_648 VDD VSS sg13g2_FILL8
XSTDFILL102_656 VDD VSS sg13g2_FILL8
XSTDFILL102_664 VDD VSS sg13g2_FILL8
XSTDFILL102_672 VDD VSS sg13g2_FILL8
XSTDFILL102_680 VDD VSS sg13g2_FILL8
XSTDFILL102_688 VDD VSS sg13g2_FILL8
XSTDFILL102_696 VDD VSS sg13g2_FILL8
XSTDFILL102_704 VDD VSS sg13g2_FILL8
XSTDFILL102_712 VDD VSS sg13g2_FILL8
XSTDFILL102_720 VDD VSS sg13g2_FILL8
XSTDFILL102_728 VDD VSS sg13g2_FILL8
XSTDFILL102_736 VDD VSS sg13g2_FILL8
XSTDFILL102_744 VDD VSS sg13g2_FILL8
XSTDFILL102_752 VDD VSS sg13g2_FILL8
XSTDFILL102_760 VDD VSS sg13g2_FILL8
XSTDFILL102_768 VDD VSS sg13g2_FILL8
XSTDFILL102_776 VDD VSS sg13g2_FILL8
XSTDFILL102_784 VDD VSS sg13g2_FILL8
XSTDFILL102_792 VDD VSS sg13g2_FILL8
XSTDFILL102_800 VDD VSS sg13g2_FILL8
XSTDFILL102_808 VDD VSS sg13g2_FILL8
XSTDFILL102_816 VDD VSS sg13g2_FILL8
XSTDFILL102_824 VDD VSS sg13g2_FILL8
XSTDFILL102_832 VDD VSS sg13g2_FILL8
XSTDFILL102_840 VDD VSS sg13g2_FILL8
XSTDFILL102_848 VDD VSS sg13g2_FILL8
XSTDFILL102_856 VDD VSS sg13g2_FILL8
XSTDFILL102_864 VDD VSS sg13g2_FILL8
XSTDFILL102_872 VDD VSS sg13g2_FILL8
XSTDFILL102_880 VDD VSS sg13g2_FILL8
XSTDFILL102_888 VDD VSS sg13g2_FILL8
XSTDFILL102_896 VDD VSS sg13g2_FILL8
XSTDFILL102_904 VDD VSS sg13g2_FILL8
XSTDFILL102_912 VDD VSS sg13g2_FILL8
XSTDFILL102_920 VDD VSS sg13g2_FILL8
XSTDFILL102_928 VDD VSS sg13g2_FILL8
XSTDFILL102_936 VDD VSS sg13g2_FILL8
XSTDFILL102_944 VDD VSS sg13g2_FILL8
XSTDFILL102_952 VDD VSS sg13g2_FILL8
XSTDFILL102_960 VDD VSS sg13g2_FILL8
XSTDFILL102_968 VDD VSS sg13g2_FILL8
XSTDFILL102_976 VDD VSS sg13g2_FILL8
XSTDFILL102_984 VDD VSS sg13g2_FILL8
XSTDFILL102_992 VDD VSS sg13g2_FILL8
XSTDFILL102_1000 VDD VSS sg13g2_FILL8
XSTDFILL102_1008 VDD VSS sg13g2_FILL8
XSTDFILL102_1016 VDD VSS sg13g2_FILL8
XSTDFILL102_1024 VDD VSS sg13g2_FILL8
XSTDFILL102_1032 VDD VSS sg13g2_FILL8
XSTDFILL102_1040 VDD VSS sg13g2_FILL8
XSTDFILL102_1048 VDD VSS sg13g2_FILL8
XSTDFILL102_1056 VDD VSS sg13g2_FILL8
XSTDFILL102_1064 VDD VSS sg13g2_FILL8
XSTDFILL102_1072 VDD VSS sg13g2_FILL8
XSTDFILL102_1080 VDD VSS sg13g2_FILL8
XSTDFILL102_1088 VDD VSS sg13g2_FILL8
XSTDFILL102_1096 VDD VSS sg13g2_FILL8
XSTDFILL102_1104 VDD VSS sg13g2_FILL8
XSTDFILL102_1112 VDD VSS sg13g2_FILL8
XSTDFILL102_1120 VDD VSS sg13g2_FILL8
XSTDFILL102_1128 VDD VSS sg13g2_FILL8
XSTDFILL102_1136 VDD VSS sg13g2_FILL8
XSTDFILL102_1144 VDD VSS sg13g2_FILL8
XSTDFILL102_1152 VDD VSS sg13g2_FILL8
XSTDFILL102_1160 VDD VSS sg13g2_FILL8
XSTDFILL102_1168 VDD VSS sg13g2_FILL8
XSTDFILL102_1176 VDD VSS sg13g2_FILL8
XSTDFILL102_1184 VDD VSS sg13g2_FILL8
XSTDFILL102_1192 VDD VSS sg13g2_FILL8
XSTDFILL102_1200 VDD VSS sg13g2_FILL8
XSTDFILL102_1208 VDD VSS sg13g2_FILL8
XSTDFILL102_1216 VDD VSS sg13g2_FILL8
XSTDFILL102_1224 VDD VSS sg13g2_FILL8
XSTDFILL102_1232 VDD VSS sg13g2_FILL8
XSTDFILL102_1240 VDD VSS sg13g2_FILL8
XSTDFILL102_1248 VDD VSS sg13g2_FILL8
XSTDFILL102_1256 VDD VSS sg13g2_FILL8
XSTDFILL102_1264 VDD VSS sg13g2_FILL8
XSTDFILL102_1272 VDD VSS sg13g2_FILL8
XSTDFILL102_1280 VDD VSS sg13g2_FILL8
XSTDFILL102_1288 VDD VSS sg13g2_FILL8
XSTDFILL102_1296 VDD VSS sg13g2_FILL8
XSTDFILL102_1304 VDD VSS sg13g2_FILL8
XSTDFILL102_1312 VDD VSS sg13g2_FILL8
XSTDFILL102_1320 VDD VSS sg13g2_FILL8
XSTDFILL102_1328 VDD VSS sg13g2_FILL8
XSTDFILL102_1336 VDD VSS sg13g2_FILL8
XSTDFILL102_1344 VDD VSS sg13g2_FILL8
XSTDFILL102_1352 VDD VSS sg13g2_FILL8
XSTDFILL102_1360 VDD VSS sg13g2_FILL8
XSTDFILL102_1368 VDD VSS sg13g2_FILL8
XSTDFILL102_1376 VDD VSS sg13g2_FILL8
XSTDFILL102_1384 VDD VSS sg13g2_FILL8
XSTDFILL102_1392 VDD VSS sg13g2_FILL8
XSTDFILL102_1400 VDD VSS sg13g2_FILL8
XSTDFILL102_1408 VDD VSS sg13g2_FILL8
XSTDFILL102_1416 VDD VSS sg13g2_FILL8
XSTDFILL102_1424 VDD VSS sg13g2_FILL8
XSTDFILL102_1432 VDD VSS sg13g2_FILL8
XSTDFILL102_1440 VDD VSS sg13g2_FILL8
XSTDFILL102_1448 VDD VSS sg13g2_FILL8
XSTDFILL102_1456 VDD VSS sg13g2_FILL8
XSTDFILL102_1464 VDD VSS sg13g2_FILL8
XSTDFILL102_1472 VDD VSS sg13g2_FILL8
XSTDFILL102_1480 VDD VSS sg13g2_FILL8
XSTDFILL102_1488 VDD VSS sg13g2_FILL8
XSTDFILL102_1496 VDD VSS sg13g2_FILL8
XSTDFILL102_1504 VDD VSS sg13g2_FILL8
XSTDFILL102_1512 VDD VSS sg13g2_FILL8
XSTDFILL102_1520 VDD VSS sg13g2_FILL8
XSTDFILL102_1528 VDD VSS sg13g2_FILL2
XSTDFILL102_1530 VDD VSS sg13g2_FILL1
XSTDFILL103_0 VDD VSS sg13g2_FILL8
XSTDFILL103_8 VDD VSS sg13g2_FILL8
XSTDFILL103_16 VDD VSS sg13g2_FILL8
XSTDFILL103_24 VDD VSS sg13g2_FILL8
XSTDFILL103_32 VDD VSS sg13g2_FILL8
XSTDFILL103_40 VDD VSS sg13g2_FILL8
XSTDFILL103_48 VDD VSS sg13g2_FILL8
XSTDFILL103_56 VDD VSS sg13g2_FILL8
XSTDFILL103_64 VDD VSS sg13g2_FILL8
XSTDFILL103_72 VDD VSS sg13g2_FILL8
XSTDFILL103_80 VDD VSS sg13g2_FILL8
XSTDFILL103_88 VDD VSS sg13g2_FILL8
XSTDFILL103_96 VDD VSS sg13g2_FILL8
XSTDFILL103_104 VDD VSS sg13g2_FILL8
XSTDFILL103_112 VDD VSS sg13g2_FILL8
XSTDFILL103_120 VDD VSS sg13g2_FILL8
XSTDFILL103_128 VDD VSS sg13g2_FILL8
XSTDFILL103_136 VDD VSS sg13g2_FILL8
XSTDFILL103_144 VDD VSS sg13g2_FILL8
XSTDFILL103_152 VDD VSS sg13g2_FILL8
XSTDFILL103_160 VDD VSS sg13g2_FILL8
XSTDFILL103_168 VDD VSS sg13g2_FILL8
XSTDFILL103_176 VDD VSS sg13g2_FILL8
XSTDFILL103_184 VDD VSS sg13g2_FILL8
XSTDFILL103_192 VDD VSS sg13g2_FILL8
XSTDFILL103_200 VDD VSS sg13g2_FILL8
XSTDFILL103_208 VDD VSS sg13g2_FILL8
XSTDFILL103_216 VDD VSS sg13g2_FILL8
XSTDFILL103_224 VDD VSS sg13g2_FILL8
XSTDFILL103_232 VDD VSS sg13g2_FILL8
XSTDFILL103_240 VDD VSS sg13g2_FILL8
XSTDFILL103_248 VDD VSS sg13g2_FILL8
XSTDFILL103_256 VDD VSS sg13g2_FILL8
XSTDFILL103_264 VDD VSS sg13g2_FILL8
XSTDFILL103_272 VDD VSS sg13g2_FILL8
XSTDFILL103_280 VDD VSS sg13g2_FILL8
XSTDFILL103_288 VDD VSS sg13g2_FILL8
XSTDFILL103_296 VDD VSS sg13g2_FILL8
XSTDFILL103_304 VDD VSS sg13g2_FILL8
XSTDFILL103_312 VDD VSS sg13g2_FILL8
XSTDFILL103_320 VDD VSS sg13g2_FILL8
XSTDFILL103_328 VDD VSS sg13g2_FILL8
XSTDFILL103_336 VDD VSS sg13g2_FILL8
XSTDFILL103_344 VDD VSS sg13g2_FILL8
XSTDFILL103_352 VDD VSS sg13g2_FILL8
XSTDFILL103_360 VDD VSS sg13g2_FILL8
XSTDFILL103_368 VDD VSS sg13g2_FILL8
XSTDFILL103_376 VDD VSS sg13g2_FILL8
XSTDFILL103_384 VDD VSS sg13g2_FILL8
XSTDFILL103_392 VDD VSS sg13g2_FILL8
XSTDFILL103_400 VDD VSS sg13g2_FILL8
XSTDFILL103_408 VDD VSS sg13g2_FILL8
XSTDFILL103_416 VDD VSS sg13g2_FILL8
XSTDFILL103_424 VDD VSS sg13g2_FILL8
XSTDFILL103_432 VDD VSS sg13g2_FILL8
XSTDFILL103_440 VDD VSS sg13g2_FILL8
XSTDFILL103_448 VDD VSS sg13g2_FILL8
XSTDFILL103_456 VDD VSS sg13g2_FILL8
XSTDFILL103_464 VDD VSS sg13g2_FILL8
XSTDFILL103_472 VDD VSS sg13g2_FILL8
XSTDFILL103_480 VDD VSS sg13g2_FILL8
XSTDFILL103_488 VDD VSS sg13g2_FILL8
XSTDFILL103_496 VDD VSS sg13g2_FILL8
XSTDFILL103_504 VDD VSS sg13g2_FILL8
XSTDFILL103_512 VDD VSS sg13g2_FILL8
XSTDFILL103_520 VDD VSS sg13g2_FILL8
XSTDFILL103_528 VDD VSS sg13g2_FILL8
XSTDFILL103_536 VDD VSS sg13g2_FILL8
XSTDFILL103_544 VDD VSS sg13g2_FILL8
XSTDFILL103_552 VDD VSS sg13g2_FILL8
XSTDFILL103_560 VDD VSS sg13g2_FILL8
XSTDFILL103_568 VDD VSS sg13g2_FILL8
XSTDFILL103_576 VDD VSS sg13g2_FILL8
XSTDFILL103_584 VDD VSS sg13g2_FILL8
XSTDFILL103_592 VDD VSS sg13g2_FILL8
XSTDFILL103_600 VDD VSS sg13g2_FILL8
XSTDFILL103_608 VDD VSS sg13g2_FILL8
XSTDFILL103_616 VDD VSS sg13g2_FILL8
XSTDFILL103_624 VDD VSS sg13g2_FILL8
XSTDFILL103_632 VDD VSS sg13g2_FILL8
XSTDFILL103_640 VDD VSS sg13g2_FILL8
XSTDFILL103_648 VDD VSS sg13g2_FILL8
XSTDFILL103_656 VDD VSS sg13g2_FILL8
XSTDFILL103_664 VDD VSS sg13g2_FILL8
XSTDFILL103_672 VDD VSS sg13g2_FILL8
XSTDFILL103_680 VDD VSS sg13g2_FILL8
XSTDFILL103_688 VDD VSS sg13g2_FILL8
XSTDFILL103_696 VDD VSS sg13g2_FILL8
XSTDFILL103_704 VDD VSS sg13g2_FILL8
XSTDFILL103_712 VDD VSS sg13g2_FILL8
XSTDFILL103_720 VDD VSS sg13g2_FILL8
XSTDFILL103_728 VDD VSS sg13g2_FILL8
XSTDFILL103_736 VDD VSS sg13g2_FILL8
XSTDFILL103_744 VDD VSS sg13g2_FILL8
XSTDFILL103_752 VDD VSS sg13g2_FILL8
XSTDFILL103_760 VDD VSS sg13g2_FILL8
XSTDFILL103_768 VDD VSS sg13g2_FILL8
XSTDFILL103_776 VDD VSS sg13g2_FILL8
XSTDFILL103_784 VDD VSS sg13g2_FILL8
XSTDFILL103_792 VDD VSS sg13g2_FILL8
XSTDFILL103_800 VDD VSS sg13g2_FILL8
XSTDFILL103_808 VDD VSS sg13g2_FILL8
XSTDFILL103_816 VDD VSS sg13g2_FILL8
XSTDFILL103_824 VDD VSS sg13g2_FILL8
XSTDFILL103_832 VDD VSS sg13g2_FILL8
XSTDFILL103_840 VDD VSS sg13g2_FILL8
XSTDFILL103_848 VDD VSS sg13g2_FILL8
XSTDFILL103_856 VDD VSS sg13g2_FILL8
XSTDFILL103_864 VDD VSS sg13g2_FILL8
XSTDFILL103_872 VDD VSS sg13g2_FILL8
XSTDFILL103_880 VDD VSS sg13g2_FILL8
XSTDFILL103_888 VDD VSS sg13g2_FILL8
XSTDFILL103_896 VDD VSS sg13g2_FILL8
XSTDFILL103_904 VDD VSS sg13g2_FILL8
XSTDFILL103_912 VDD VSS sg13g2_FILL8
XSTDFILL103_920 VDD VSS sg13g2_FILL8
XSTDFILL103_928 VDD VSS sg13g2_FILL8
XSTDFILL103_936 VDD VSS sg13g2_FILL8
XSTDFILL103_944 VDD VSS sg13g2_FILL8
XSTDFILL103_952 VDD VSS sg13g2_FILL8
XSTDFILL103_960 VDD VSS sg13g2_FILL8
XSTDFILL103_968 VDD VSS sg13g2_FILL8
XSTDFILL103_976 VDD VSS sg13g2_FILL8
XSTDFILL103_984 VDD VSS sg13g2_FILL8
XSTDFILL103_992 VDD VSS sg13g2_FILL8
XSTDFILL103_1000 VDD VSS sg13g2_FILL8
XSTDFILL103_1008 VDD VSS sg13g2_FILL8
XSTDFILL103_1016 VDD VSS sg13g2_FILL8
XSTDFILL103_1024 VDD VSS sg13g2_FILL8
XSTDFILL103_1032 VDD VSS sg13g2_FILL8
XSTDFILL103_1040 VDD VSS sg13g2_FILL8
XSTDFILL103_1048 VDD VSS sg13g2_FILL8
XSTDFILL103_1056 VDD VSS sg13g2_FILL8
XSTDFILL103_1064 VDD VSS sg13g2_FILL8
XSTDFILL103_1072 VDD VSS sg13g2_FILL8
XSTDFILL103_1080 VDD VSS sg13g2_FILL8
XSTDFILL103_1088 VDD VSS sg13g2_FILL8
XSTDFILL103_1096 VDD VSS sg13g2_FILL8
XSTDFILL103_1104 VDD VSS sg13g2_FILL8
XSTDFILL103_1112 VDD VSS sg13g2_FILL8
XSTDFILL103_1120 VDD VSS sg13g2_FILL8
XSTDFILL103_1128 VDD VSS sg13g2_FILL8
XSTDFILL103_1136 VDD VSS sg13g2_FILL8
XSTDFILL103_1144 VDD VSS sg13g2_FILL8
XSTDFILL103_1152 VDD VSS sg13g2_FILL8
XSTDFILL103_1160 VDD VSS sg13g2_FILL8
XSTDFILL103_1168 VDD VSS sg13g2_FILL8
XSTDFILL103_1176 VDD VSS sg13g2_FILL8
XSTDFILL103_1184 VDD VSS sg13g2_FILL8
XSTDFILL103_1192 VDD VSS sg13g2_FILL8
XSTDFILL103_1200 VDD VSS sg13g2_FILL8
XSTDFILL103_1208 VDD VSS sg13g2_FILL8
XSTDFILL103_1216 VDD VSS sg13g2_FILL8
XSTDFILL103_1224 VDD VSS sg13g2_FILL8
XSTDFILL103_1232 VDD VSS sg13g2_FILL8
XSTDFILL103_1240 VDD VSS sg13g2_FILL8
XSTDFILL103_1248 VDD VSS sg13g2_FILL8
XSTDFILL103_1256 VDD VSS sg13g2_FILL8
XSTDFILL103_1264 VDD VSS sg13g2_FILL8
XSTDFILL103_1272 VDD VSS sg13g2_FILL8
XSTDFILL103_1280 VDD VSS sg13g2_FILL8
XSTDFILL103_1288 VDD VSS sg13g2_FILL8
XSTDFILL103_1296 VDD VSS sg13g2_FILL8
XSTDFILL103_1304 VDD VSS sg13g2_FILL8
XSTDFILL103_1312 VDD VSS sg13g2_FILL8
XSTDFILL103_1320 VDD VSS sg13g2_FILL8
XSTDFILL103_1328 VDD VSS sg13g2_FILL8
XSTDFILL103_1336 VDD VSS sg13g2_FILL8
XSTDFILL103_1344 VDD VSS sg13g2_FILL8
XSTDFILL103_1352 VDD VSS sg13g2_FILL8
XSTDFILL103_1360 VDD VSS sg13g2_FILL8
XSTDFILL103_1368 VDD VSS sg13g2_FILL8
XSTDFILL103_1376 VDD VSS sg13g2_FILL8
XSTDFILL103_1384 VDD VSS sg13g2_FILL8
XSTDFILL103_1392 VDD VSS sg13g2_FILL8
XSTDFILL103_1400 VDD VSS sg13g2_FILL8
XSTDFILL103_1408 VDD VSS sg13g2_FILL8
XSTDFILL103_1416 VDD VSS sg13g2_FILL8
XSTDFILL103_1424 VDD VSS sg13g2_FILL8
XSTDFILL103_1432 VDD VSS sg13g2_FILL8
XSTDFILL103_1440 VDD VSS sg13g2_FILL8
XSTDFILL103_1448 VDD VSS sg13g2_FILL8
XSTDFILL103_1456 VDD VSS sg13g2_FILL8
XSTDFILL103_1464 VDD VSS sg13g2_FILL8
XSTDFILL103_1472 VDD VSS sg13g2_FILL8
XSTDFILL103_1480 VDD VSS sg13g2_FILL8
XSTDFILL103_1488 VDD VSS sg13g2_FILL8
XSTDFILL103_1496 VDD VSS sg13g2_FILL8
XSTDFILL103_1504 VDD VSS sg13g2_FILL8
XSTDFILL103_1512 VDD VSS sg13g2_FILL8
XSTDFILL103_1520 VDD VSS sg13g2_FILL8
XSTDFILL103_1528 VDD VSS sg13g2_FILL2
XSTDFILL103_1530 VDD VSS sg13g2_FILL1
XSTDFILL104_0 VDD VSS sg13g2_FILL8
XSTDFILL104_8 VDD VSS sg13g2_FILL8
XSTDFILL104_16 VDD VSS sg13g2_FILL8
XSTDFILL104_24 VDD VSS sg13g2_FILL8
XSTDFILL104_32 VDD VSS sg13g2_FILL8
XSTDFILL104_40 VDD VSS sg13g2_FILL8
XSTDFILL104_48 VDD VSS sg13g2_FILL8
XSTDFILL104_56 VDD VSS sg13g2_FILL8
XSTDFILL104_64 VDD VSS sg13g2_FILL8
XSTDFILL104_72 VDD VSS sg13g2_FILL8
XSTDFILL104_80 VDD VSS sg13g2_FILL8
XSTDFILL104_88 VDD VSS sg13g2_FILL8
XSTDFILL104_96 VDD VSS sg13g2_FILL8
XSTDFILL104_104 VDD VSS sg13g2_FILL8
XSTDFILL104_112 VDD VSS sg13g2_FILL8
XSTDFILL104_120 VDD VSS sg13g2_FILL8
XSTDFILL104_128 VDD VSS sg13g2_FILL8
XSTDFILL104_136 VDD VSS sg13g2_FILL8
XSTDFILL104_144 VDD VSS sg13g2_FILL8
XSTDFILL104_152 VDD VSS sg13g2_FILL8
XSTDFILL104_160 VDD VSS sg13g2_FILL8
XSTDFILL104_168 VDD VSS sg13g2_FILL8
XSTDFILL104_176 VDD VSS sg13g2_FILL8
XSTDFILL104_184 VDD VSS sg13g2_FILL8
XSTDFILL104_192 VDD VSS sg13g2_FILL8
XSTDFILL104_200 VDD VSS sg13g2_FILL8
XSTDFILL104_208 VDD VSS sg13g2_FILL8
XSTDFILL104_216 VDD VSS sg13g2_FILL8
XSTDFILL104_224 VDD VSS sg13g2_FILL8
XSTDFILL104_232 VDD VSS sg13g2_FILL8
XSTDFILL104_240 VDD VSS sg13g2_FILL8
XSTDFILL104_248 VDD VSS sg13g2_FILL8
XSTDFILL104_256 VDD VSS sg13g2_FILL8
XSTDFILL104_264 VDD VSS sg13g2_FILL8
XSTDFILL104_272 VDD VSS sg13g2_FILL8
XSTDFILL104_280 VDD VSS sg13g2_FILL8
XSTDFILL104_288 VDD VSS sg13g2_FILL8
XSTDFILL104_296 VDD VSS sg13g2_FILL8
XSTDFILL104_304 VDD VSS sg13g2_FILL8
XSTDFILL104_312 VDD VSS sg13g2_FILL8
XSTDFILL104_320 VDD VSS sg13g2_FILL8
XSTDFILL104_328 VDD VSS sg13g2_FILL8
XSTDFILL104_336 VDD VSS sg13g2_FILL8
XSTDFILL104_344 VDD VSS sg13g2_FILL8
XSTDFILL104_352 VDD VSS sg13g2_FILL8
XSTDFILL104_360 VDD VSS sg13g2_FILL8
XSTDFILL104_368 VDD VSS sg13g2_FILL8
XSTDFILL104_376 VDD VSS sg13g2_FILL8
XSTDFILL104_384 VDD VSS sg13g2_FILL8
XSTDFILL104_392 VDD VSS sg13g2_FILL8
XSTDFILL104_400 VDD VSS sg13g2_FILL8
XSTDFILL104_408 VDD VSS sg13g2_FILL8
XSTDFILL104_416 VDD VSS sg13g2_FILL8
XSTDFILL104_424 VDD VSS sg13g2_FILL8
XSTDFILL104_432 VDD VSS sg13g2_FILL8
XSTDFILL104_440 VDD VSS sg13g2_FILL8
XSTDFILL104_448 VDD VSS sg13g2_FILL8
XSTDFILL104_456 VDD VSS sg13g2_FILL8
XSTDFILL104_464 VDD VSS sg13g2_FILL8
XSTDFILL104_472 VDD VSS sg13g2_FILL8
XSTDFILL104_480 VDD VSS sg13g2_FILL8
XSTDFILL104_488 VDD VSS sg13g2_FILL8
XSTDFILL104_496 VDD VSS sg13g2_FILL8
XSTDFILL104_504 VDD VSS sg13g2_FILL8
XSTDFILL104_512 VDD VSS sg13g2_FILL8
XSTDFILL104_520 VDD VSS sg13g2_FILL8
XSTDFILL104_528 VDD VSS sg13g2_FILL8
XSTDFILL104_536 VDD VSS sg13g2_FILL8
XSTDFILL104_544 VDD VSS sg13g2_FILL8
XSTDFILL104_552 VDD VSS sg13g2_FILL8
XSTDFILL104_560 VDD VSS sg13g2_FILL8
XSTDFILL104_568 VDD VSS sg13g2_FILL8
XSTDFILL104_576 VDD VSS sg13g2_FILL8
XSTDFILL104_584 VDD VSS sg13g2_FILL8
XSTDFILL104_592 VDD VSS sg13g2_FILL8
XSTDFILL104_600 VDD VSS sg13g2_FILL8
XSTDFILL104_608 VDD VSS sg13g2_FILL8
XSTDFILL104_616 VDD VSS sg13g2_FILL8
XSTDFILL104_624 VDD VSS sg13g2_FILL8
XSTDFILL104_632 VDD VSS sg13g2_FILL8
XSTDFILL104_640 VDD VSS sg13g2_FILL8
XSTDFILL104_648 VDD VSS sg13g2_FILL8
XSTDFILL104_656 VDD VSS sg13g2_FILL8
XSTDFILL104_664 VDD VSS sg13g2_FILL8
XSTDFILL104_672 VDD VSS sg13g2_FILL8
XSTDFILL104_680 VDD VSS sg13g2_FILL8
XSTDFILL104_688 VDD VSS sg13g2_FILL8
XSTDFILL104_696 VDD VSS sg13g2_FILL8
XSTDFILL104_704 VDD VSS sg13g2_FILL8
XSTDFILL104_712 VDD VSS sg13g2_FILL8
XSTDFILL104_720 VDD VSS sg13g2_FILL8
XSTDFILL104_728 VDD VSS sg13g2_FILL8
XSTDFILL104_736 VDD VSS sg13g2_FILL8
XSTDFILL104_744 VDD VSS sg13g2_FILL8
XSTDFILL104_752 VDD VSS sg13g2_FILL8
XSTDFILL104_760 VDD VSS sg13g2_FILL8
XSTDFILL104_768 VDD VSS sg13g2_FILL8
XSTDFILL104_776 VDD VSS sg13g2_FILL8
XSTDFILL104_784 VDD VSS sg13g2_FILL8
XSTDFILL104_792 VDD VSS sg13g2_FILL8
XSTDFILL104_800 VDD VSS sg13g2_FILL8
XSTDFILL104_808 VDD VSS sg13g2_FILL8
XSTDFILL104_816 VDD VSS sg13g2_FILL8
XSTDFILL104_824 VDD VSS sg13g2_FILL8
XSTDFILL104_832 VDD VSS sg13g2_FILL8
XSTDFILL104_840 VDD VSS sg13g2_FILL8
XSTDFILL104_848 VDD VSS sg13g2_FILL8
XSTDFILL104_856 VDD VSS sg13g2_FILL8
XSTDFILL104_864 VDD VSS sg13g2_FILL8
XSTDFILL104_872 VDD VSS sg13g2_FILL8
XSTDFILL104_880 VDD VSS sg13g2_FILL8
XSTDFILL104_888 VDD VSS sg13g2_FILL8
XSTDFILL104_896 VDD VSS sg13g2_FILL8
XSTDFILL104_904 VDD VSS sg13g2_FILL8
XSTDFILL104_912 VDD VSS sg13g2_FILL8
XSTDFILL104_920 VDD VSS sg13g2_FILL8
XSTDFILL104_928 VDD VSS sg13g2_FILL8
XSTDFILL104_936 VDD VSS sg13g2_FILL8
XSTDFILL104_944 VDD VSS sg13g2_FILL8
XSTDFILL104_952 VDD VSS sg13g2_FILL8
XSTDFILL104_960 VDD VSS sg13g2_FILL8
XSTDFILL104_968 VDD VSS sg13g2_FILL8
XSTDFILL104_976 VDD VSS sg13g2_FILL8
XSTDFILL104_984 VDD VSS sg13g2_FILL8
XSTDFILL104_992 VDD VSS sg13g2_FILL8
XSTDFILL104_1000 VDD VSS sg13g2_FILL8
XSTDFILL104_1008 VDD VSS sg13g2_FILL8
XSTDFILL104_1016 VDD VSS sg13g2_FILL8
XSTDFILL104_1024 VDD VSS sg13g2_FILL8
XSTDFILL104_1032 VDD VSS sg13g2_FILL8
XSTDFILL104_1040 VDD VSS sg13g2_FILL8
XSTDFILL104_1048 VDD VSS sg13g2_FILL8
XSTDFILL104_1056 VDD VSS sg13g2_FILL8
XSTDFILL104_1064 VDD VSS sg13g2_FILL8
XSTDFILL104_1072 VDD VSS sg13g2_FILL8
XSTDFILL104_1080 VDD VSS sg13g2_FILL8
XSTDFILL104_1088 VDD VSS sg13g2_FILL8
XSTDFILL104_1096 VDD VSS sg13g2_FILL8
XSTDFILL104_1104 VDD VSS sg13g2_FILL8
XSTDFILL104_1112 VDD VSS sg13g2_FILL8
XSTDFILL104_1120 VDD VSS sg13g2_FILL8
XSTDFILL104_1128 VDD VSS sg13g2_FILL8
XSTDFILL104_1136 VDD VSS sg13g2_FILL8
XSTDFILL104_1144 VDD VSS sg13g2_FILL8
XSTDFILL104_1152 VDD VSS sg13g2_FILL8
XSTDFILL104_1160 VDD VSS sg13g2_FILL8
XSTDFILL104_1168 VDD VSS sg13g2_FILL8
XSTDFILL104_1176 VDD VSS sg13g2_FILL8
XSTDFILL104_1184 VDD VSS sg13g2_FILL8
XSTDFILL104_1192 VDD VSS sg13g2_FILL8
XSTDFILL104_1200 VDD VSS sg13g2_FILL8
XSTDFILL104_1208 VDD VSS sg13g2_FILL8
XSTDFILL104_1216 VDD VSS sg13g2_FILL8
XSTDFILL104_1224 VDD VSS sg13g2_FILL8
XSTDFILL104_1232 VDD VSS sg13g2_FILL8
XSTDFILL104_1240 VDD VSS sg13g2_FILL8
XSTDFILL104_1248 VDD VSS sg13g2_FILL8
XSTDFILL104_1256 VDD VSS sg13g2_FILL8
XSTDFILL104_1264 VDD VSS sg13g2_FILL8
XSTDFILL104_1272 VDD VSS sg13g2_FILL8
XSTDFILL104_1280 VDD VSS sg13g2_FILL8
XSTDFILL104_1288 VDD VSS sg13g2_FILL8
XSTDFILL104_1296 VDD VSS sg13g2_FILL8
XSTDFILL104_1304 VDD VSS sg13g2_FILL8
XSTDFILL104_1312 VDD VSS sg13g2_FILL8
XSTDFILL104_1320 VDD VSS sg13g2_FILL8
XSTDFILL104_1328 VDD VSS sg13g2_FILL8
XSTDFILL104_1336 VDD VSS sg13g2_FILL8
XSTDFILL104_1344 VDD VSS sg13g2_FILL8
XSTDFILL104_1352 VDD VSS sg13g2_FILL8
XSTDFILL104_1360 VDD VSS sg13g2_FILL8
XSTDFILL104_1368 VDD VSS sg13g2_FILL8
XSTDFILL104_1376 VDD VSS sg13g2_FILL8
XSTDFILL104_1384 VDD VSS sg13g2_FILL8
XSTDFILL104_1392 VDD VSS sg13g2_FILL8
XSTDFILL104_1400 VDD VSS sg13g2_FILL8
XSTDFILL104_1408 VDD VSS sg13g2_FILL8
XSTDFILL104_1416 VDD VSS sg13g2_FILL8
XSTDFILL104_1424 VDD VSS sg13g2_FILL8
XSTDFILL104_1432 VDD VSS sg13g2_FILL8
XSTDFILL104_1440 VDD VSS sg13g2_FILL8
XSTDFILL104_1448 VDD VSS sg13g2_FILL8
XSTDFILL104_1456 VDD VSS sg13g2_FILL8
XSTDFILL104_1464 VDD VSS sg13g2_FILL8
XSTDFILL104_1472 VDD VSS sg13g2_FILL8
XSTDFILL104_1480 VDD VSS sg13g2_FILL8
XSTDFILL104_1488 VDD VSS sg13g2_FILL8
XSTDFILL104_1496 VDD VSS sg13g2_FILL8
XSTDFILL104_1504 VDD VSS sg13g2_FILL8
XSTDFILL104_1512 VDD VSS sg13g2_FILL8
XSTDFILL104_1520 VDD VSS sg13g2_FILL8
XSTDFILL104_1528 VDD VSS sg13g2_FILL2
XSTDFILL104_1530 VDD VSS sg13g2_FILL1
XSTDFILL105_0 VDD VSS sg13g2_FILL8
XSTDFILL105_8 VDD VSS sg13g2_FILL8
XSTDFILL105_16 VDD VSS sg13g2_FILL8
XSTDFILL105_24 VDD VSS sg13g2_FILL8
XSTDFILL105_32 VDD VSS sg13g2_FILL8
XSTDFILL105_40 VDD VSS sg13g2_FILL8
XSTDFILL105_48 VDD VSS sg13g2_FILL8
XSTDFILL105_56 VDD VSS sg13g2_FILL8
XSTDFILL105_64 VDD VSS sg13g2_FILL8
XSTDFILL105_72 VDD VSS sg13g2_FILL8
XSTDFILL105_80 VDD VSS sg13g2_FILL8
XSTDFILL105_88 VDD VSS sg13g2_FILL8
XSTDFILL105_96 VDD VSS sg13g2_FILL8
XSTDFILL105_104 VDD VSS sg13g2_FILL8
XSTDFILL105_112 VDD VSS sg13g2_FILL8
XSTDFILL105_120 VDD VSS sg13g2_FILL8
XSTDFILL105_128 VDD VSS sg13g2_FILL8
XSTDFILL105_136 VDD VSS sg13g2_FILL8
XSTDFILL105_144 VDD VSS sg13g2_FILL8
XSTDFILL105_152 VDD VSS sg13g2_FILL8
XSTDFILL105_160 VDD VSS sg13g2_FILL8
XSTDFILL105_168 VDD VSS sg13g2_FILL8
XSTDFILL105_176 VDD VSS sg13g2_FILL8
XSTDFILL105_184 VDD VSS sg13g2_FILL8
XSTDFILL105_192 VDD VSS sg13g2_FILL8
XSTDFILL105_200 VDD VSS sg13g2_FILL8
XSTDFILL105_208 VDD VSS sg13g2_FILL8
XSTDFILL105_216 VDD VSS sg13g2_FILL8
XSTDFILL105_224 VDD VSS sg13g2_FILL8
XSTDFILL105_232 VDD VSS sg13g2_FILL8
XSTDFILL105_240 VDD VSS sg13g2_FILL8
XSTDFILL105_248 VDD VSS sg13g2_FILL8
XSTDFILL105_256 VDD VSS sg13g2_FILL8
XSTDFILL105_264 VDD VSS sg13g2_FILL8
XSTDFILL105_272 VDD VSS sg13g2_FILL8
XSTDFILL105_280 VDD VSS sg13g2_FILL8
XSTDFILL105_288 VDD VSS sg13g2_FILL8
XSTDFILL105_296 VDD VSS sg13g2_FILL8
XSTDFILL105_304 VDD VSS sg13g2_FILL8
XSTDFILL105_312 VDD VSS sg13g2_FILL8
XSTDFILL105_320 VDD VSS sg13g2_FILL8
XSTDFILL105_328 VDD VSS sg13g2_FILL8
XSTDFILL105_336 VDD VSS sg13g2_FILL8
XSTDFILL105_344 VDD VSS sg13g2_FILL8
XSTDFILL105_352 VDD VSS sg13g2_FILL8
XSTDFILL105_360 VDD VSS sg13g2_FILL8
XSTDFILL105_368 VDD VSS sg13g2_FILL8
XSTDFILL105_376 VDD VSS sg13g2_FILL8
XSTDFILL105_384 VDD VSS sg13g2_FILL8
XSTDFILL105_392 VDD VSS sg13g2_FILL8
XSTDFILL105_400 VDD VSS sg13g2_FILL8
XSTDFILL105_408 VDD VSS sg13g2_FILL8
XSTDFILL105_416 VDD VSS sg13g2_FILL8
XSTDFILL105_424 VDD VSS sg13g2_FILL8
XSTDFILL105_432 VDD VSS sg13g2_FILL8
XSTDFILL105_440 VDD VSS sg13g2_FILL8
XSTDFILL105_448 VDD VSS sg13g2_FILL8
XSTDFILL105_456 VDD VSS sg13g2_FILL8
XSTDFILL105_464 VDD VSS sg13g2_FILL8
XSTDFILL105_472 VDD VSS sg13g2_FILL8
XSTDFILL105_480 VDD VSS sg13g2_FILL8
XSTDFILL105_488 VDD VSS sg13g2_FILL8
XSTDFILL105_496 VDD VSS sg13g2_FILL8
XSTDFILL105_504 VDD VSS sg13g2_FILL8
XSTDFILL105_512 VDD VSS sg13g2_FILL8
XSTDFILL105_520 VDD VSS sg13g2_FILL8
XSTDFILL105_528 VDD VSS sg13g2_FILL8
XSTDFILL105_536 VDD VSS sg13g2_FILL8
XSTDFILL105_544 VDD VSS sg13g2_FILL8
XSTDFILL105_552 VDD VSS sg13g2_FILL8
XSTDFILL105_560 VDD VSS sg13g2_FILL8
XSTDFILL105_568 VDD VSS sg13g2_FILL8
XSTDFILL105_576 VDD VSS sg13g2_FILL8
XSTDFILL105_584 VDD VSS sg13g2_FILL8
XSTDFILL105_592 VDD VSS sg13g2_FILL8
XSTDFILL105_600 VDD VSS sg13g2_FILL8
XSTDFILL105_608 VDD VSS sg13g2_FILL8
XSTDFILL105_616 VDD VSS sg13g2_FILL8
XSTDFILL105_624 VDD VSS sg13g2_FILL8
XSTDFILL105_632 VDD VSS sg13g2_FILL8
XSTDFILL105_640 VDD VSS sg13g2_FILL8
XSTDFILL105_648 VDD VSS sg13g2_FILL8
XSTDFILL105_656 VDD VSS sg13g2_FILL8
XSTDFILL105_664 VDD VSS sg13g2_FILL8
XSTDFILL105_672 VDD VSS sg13g2_FILL8
XSTDFILL105_680 VDD VSS sg13g2_FILL8
XSTDFILL105_688 VDD VSS sg13g2_FILL8
XSTDFILL105_696 VDD VSS sg13g2_FILL8
XSTDFILL105_704 VDD VSS sg13g2_FILL8
XSTDFILL105_712 VDD VSS sg13g2_FILL8
XSTDFILL105_720 VDD VSS sg13g2_FILL8
XSTDFILL105_728 VDD VSS sg13g2_FILL8
XSTDFILL105_736 VDD VSS sg13g2_FILL8
XSTDFILL105_744 VDD VSS sg13g2_FILL8
XSTDFILL105_752 VDD VSS sg13g2_FILL8
XSTDFILL105_760 VDD VSS sg13g2_FILL8
XSTDFILL105_768 VDD VSS sg13g2_FILL8
XSTDFILL105_776 VDD VSS sg13g2_FILL8
XSTDFILL105_784 VDD VSS sg13g2_FILL8
XSTDFILL105_792 VDD VSS sg13g2_FILL8
XSTDFILL105_800 VDD VSS sg13g2_FILL8
XSTDFILL105_808 VDD VSS sg13g2_FILL8
XSTDFILL105_816 VDD VSS sg13g2_FILL8
XSTDFILL105_824 VDD VSS sg13g2_FILL8
XSTDFILL105_832 VDD VSS sg13g2_FILL8
XSTDFILL105_840 VDD VSS sg13g2_FILL8
XSTDFILL105_848 VDD VSS sg13g2_FILL8
XSTDFILL105_856 VDD VSS sg13g2_FILL8
XSTDFILL105_864 VDD VSS sg13g2_FILL8
XSTDFILL105_872 VDD VSS sg13g2_FILL8
XSTDFILL105_880 VDD VSS sg13g2_FILL8
XSTDFILL105_888 VDD VSS sg13g2_FILL8
XSTDFILL105_896 VDD VSS sg13g2_FILL8
XSTDFILL105_904 VDD VSS sg13g2_FILL8
XSTDFILL105_912 VDD VSS sg13g2_FILL8
XSTDFILL105_920 VDD VSS sg13g2_FILL8
XSTDFILL105_928 VDD VSS sg13g2_FILL8
XSTDFILL105_936 VDD VSS sg13g2_FILL8
XSTDFILL105_944 VDD VSS sg13g2_FILL8
XSTDFILL105_952 VDD VSS sg13g2_FILL8
XSTDFILL105_960 VDD VSS sg13g2_FILL8
XSTDFILL105_968 VDD VSS sg13g2_FILL8
XSTDFILL105_976 VDD VSS sg13g2_FILL8
XSTDFILL105_984 VDD VSS sg13g2_FILL8
XSTDFILL105_992 VDD VSS sg13g2_FILL8
XSTDFILL105_1000 VDD VSS sg13g2_FILL8
XSTDFILL105_1008 VDD VSS sg13g2_FILL8
XSTDFILL105_1016 VDD VSS sg13g2_FILL8
XSTDFILL105_1024 VDD VSS sg13g2_FILL8
XSTDFILL105_1032 VDD VSS sg13g2_FILL8
XSTDFILL105_1040 VDD VSS sg13g2_FILL8
XSTDFILL105_1048 VDD VSS sg13g2_FILL8
XSTDFILL105_1056 VDD VSS sg13g2_FILL8
XSTDFILL105_1064 VDD VSS sg13g2_FILL8
XSTDFILL105_1072 VDD VSS sg13g2_FILL8
XSTDFILL105_1080 VDD VSS sg13g2_FILL8
XSTDFILL105_1088 VDD VSS sg13g2_FILL8
XSTDFILL105_1096 VDD VSS sg13g2_FILL8
XSTDFILL105_1104 VDD VSS sg13g2_FILL8
XSTDFILL105_1112 VDD VSS sg13g2_FILL8
XSTDFILL105_1120 VDD VSS sg13g2_FILL8
XSTDFILL105_1128 VDD VSS sg13g2_FILL8
XSTDFILL105_1136 VDD VSS sg13g2_FILL8
XSTDFILL105_1144 VDD VSS sg13g2_FILL8
XSTDFILL105_1152 VDD VSS sg13g2_FILL8
XSTDFILL105_1160 VDD VSS sg13g2_FILL8
XSTDFILL105_1168 VDD VSS sg13g2_FILL8
XSTDFILL105_1176 VDD VSS sg13g2_FILL8
XSTDFILL105_1184 VDD VSS sg13g2_FILL8
XSTDFILL105_1192 VDD VSS sg13g2_FILL8
XSTDFILL105_1200 VDD VSS sg13g2_FILL8
XSTDFILL105_1208 VDD VSS sg13g2_FILL8
XSTDFILL105_1216 VDD VSS sg13g2_FILL8
XSTDFILL105_1224 VDD VSS sg13g2_FILL8
XSTDFILL105_1232 VDD VSS sg13g2_FILL8
XSTDFILL105_1240 VDD VSS sg13g2_FILL8
XSTDFILL105_1248 VDD VSS sg13g2_FILL8
XSTDFILL105_1256 VDD VSS sg13g2_FILL8
XSTDFILL105_1264 VDD VSS sg13g2_FILL8
XSTDFILL105_1272 VDD VSS sg13g2_FILL8
XSTDFILL105_1280 VDD VSS sg13g2_FILL8
XSTDFILL105_1288 VDD VSS sg13g2_FILL8
XSTDFILL105_1296 VDD VSS sg13g2_FILL8
XSTDFILL105_1304 VDD VSS sg13g2_FILL8
XSTDFILL105_1312 VDD VSS sg13g2_FILL8
XSTDFILL105_1320 VDD VSS sg13g2_FILL8
XSTDFILL105_1328 VDD VSS sg13g2_FILL8
XSTDFILL105_1336 VDD VSS sg13g2_FILL8
XSTDFILL105_1344 VDD VSS sg13g2_FILL8
XSTDFILL105_1352 VDD VSS sg13g2_FILL8
XSTDFILL105_1360 VDD VSS sg13g2_FILL8
XSTDFILL105_1368 VDD VSS sg13g2_FILL8
XSTDFILL105_1376 VDD VSS sg13g2_FILL8
XSTDFILL105_1384 VDD VSS sg13g2_FILL8
XSTDFILL105_1392 VDD VSS sg13g2_FILL8
XSTDFILL105_1400 VDD VSS sg13g2_FILL8
XSTDFILL105_1408 VDD VSS sg13g2_FILL8
XSTDFILL105_1416 VDD VSS sg13g2_FILL8
XSTDFILL105_1424 VDD VSS sg13g2_FILL8
XSTDFILL105_1432 VDD VSS sg13g2_FILL8
XSTDFILL105_1440 VDD VSS sg13g2_FILL8
XSTDFILL105_1448 VDD VSS sg13g2_FILL8
XSTDFILL105_1456 VDD VSS sg13g2_FILL8
XSTDFILL105_1464 VDD VSS sg13g2_FILL8
XSTDFILL105_1472 VDD VSS sg13g2_FILL8
XSTDFILL105_1480 VDD VSS sg13g2_FILL8
XSTDFILL105_1488 VDD VSS sg13g2_FILL8
XSTDFILL105_1496 VDD VSS sg13g2_FILL8
XSTDFILL105_1504 VDD VSS sg13g2_FILL8
XSTDFILL105_1512 VDD VSS sg13g2_FILL8
XSTDFILL105_1520 VDD VSS sg13g2_FILL8
XSTDFILL105_1528 VDD VSS sg13g2_FILL2
XSTDFILL105_1530 VDD VSS sg13g2_FILL1
XSTDFILL106_0 VDD VSS sg13g2_FILL8
XSTDFILL106_8 VDD VSS sg13g2_FILL8
XSTDFILL106_16 VDD VSS sg13g2_FILL8
XSTDFILL106_24 VDD VSS sg13g2_FILL8
XSTDFILL106_32 VDD VSS sg13g2_FILL8
XSTDFILL106_40 VDD VSS sg13g2_FILL8
XSTDFILL106_48 VDD VSS sg13g2_FILL8
XSTDFILL106_56 VDD VSS sg13g2_FILL8
XSTDFILL106_64 VDD VSS sg13g2_FILL8
XSTDFILL106_72 VDD VSS sg13g2_FILL8
XSTDFILL106_80 VDD VSS sg13g2_FILL8
XSTDFILL106_88 VDD VSS sg13g2_FILL8
XSTDFILL106_96 VDD VSS sg13g2_FILL8
XSTDFILL106_104 VDD VSS sg13g2_FILL8
XSTDFILL106_112 VDD VSS sg13g2_FILL8
XSTDFILL106_120 VDD VSS sg13g2_FILL8
XSTDFILL106_128 VDD VSS sg13g2_FILL8
XSTDFILL106_136 VDD VSS sg13g2_FILL8
XSTDFILL106_144 VDD VSS sg13g2_FILL8
XSTDFILL106_152 VDD VSS sg13g2_FILL8
XSTDFILL106_160 VDD VSS sg13g2_FILL8
XSTDFILL106_168 VDD VSS sg13g2_FILL8
XSTDFILL106_176 VDD VSS sg13g2_FILL8
XSTDFILL106_184 VDD VSS sg13g2_FILL8
XSTDFILL106_192 VDD VSS sg13g2_FILL8
XSTDFILL106_200 VDD VSS sg13g2_FILL8
XSTDFILL106_208 VDD VSS sg13g2_FILL8
XSTDFILL106_216 VDD VSS sg13g2_FILL8
XSTDFILL106_224 VDD VSS sg13g2_FILL8
XSTDFILL106_232 VDD VSS sg13g2_FILL8
XSTDFILL106_240 VDD VSS sg13g2_FILL8
XSTDFILL106_248 VDD VSS sg13g2_FILL8
XSTDFILL106_256 VDD VSS sg13g2_FILL8
XSTDFILL106_264 VDD VSS sg13g2_FILL8
XSTDFILL106_272 VDD VSS sg13g2_FILL8
XSTDFILL106_280 VDD VSS sg13g2_FILL8
XSTDFILL106_288 VDD VSS sg13g2_FILL8
XSTDFILL106_296 VDD VSS sg13g2_FILL8
XSTDFILL106_304 VDD VSS sg13g2_FILL8
XSTDFILL106_312 VDD VSS sg13g2_FILL8
XSTDFILL106_320 VDD VSS sg13g2_FILL8
XSTDFILL106_328 VDD VSS sg13g2_FILL8
XSTDFILL106_336 VDD VSS sg13g2_FILL8
XSTDFILL106_344 VDD VSS sg13g2_FILL8
XSTDFILL106_352 VDD VSS sg13g2_FILL8
XSTDFILL106_360 VDD VSS sg13g2_FILL8
XSTDFILL106_368 VDD VSS sg13g2_FILL8
XSTDFILL106_376 VDD VSS sg13g2_FILL8
XSTDFILL106_384 VDD VSS sg13g2_FILL8
XSTDFILL106_392 VDD VSS sg13g2_FILL8
XSTDFILL106_400 VDD VSS sg13g2_FILL8
XSTDFILL106_408 VDD VSS sg13g2_FILL8
XSTDFILL106_416 VDD VSS sg13g2_FILL8
XSTDFILL106_424 VDD VSS sg13g2_FILL8
XSTDFILL106_432 VDD VSS sg13g2_FILL8
XSTDFILL106_440 VDD VSS sg13g2_FILL8
XSTDFILL106_448 VDD VSS sg13g2_FILL8
XSTDFILL106_456 VDD VSS sg13g2_FILL8
XSTDFILL106_464 VDD VSS sg13g2_FILL8
XSTDFILL106_472 VDD VSS sg13g2_FILL8
XSTDFILL106_480 VDD VSS sg13g2_FILL8
XSTDFILL106_488 VDD VSS sg13g2_FILL8
XSTDFILL106_496 VDD VSS sg13g2_FILL8
XSTDFILL106_504 VDD VSS sg13g2_FILL8
XSTDFILL106_512 VDD VSS sg13g2_FILL8
XSTDFILL106_520 VDD VSS sg13g2_FILL8
XSTDFILL106_528 VDD VSS sg13g2_FILL8
XSTDFILL106_536 VDD VSS sg13g2_FILL8
XSTDFILL106_544 VDD VSS sg13g2_FILL8
XSTDFILL106_552 VDD VSS sg13g2_FILL8
XSTDFILL106_560 VDD VSS sg13g2_FILL8
XSTDFILL106_568 VDD VSS sg13g2_FILL8
XSTDFILL106_576 VDD VSS sg13g2_FILL8
XSTDFILL106_584 VDD VSS sg13g2_FILL8
XSTDFILL106_592 VDD VSS sg13g2_FILL8
XSTDFILL106_600 VDD VSS sg13g2_FILL8
XSTDFILL106_608 VDD VSS sg13g2_FILL8
XSTDFILL106_616 VDD VSS sg13g2_FILL8
XSTDFILL106_624 VDD VSS sg13g2_FILL8
XSTDFILL106_632 VDD VSS sg13g2_FILL8
XSTDFILL106_640 VDD VSS sg13g2_FILL8
XSTDFILL106_648 VDD VSS sg13g2_FILL8
XSTDFILL106_656 VDD VSS sg13g2_FILL8
XSTDFILL106_664 VDD VSS sg13g2_FILL8
XSTDFILL106_672 VDD VSS sg13g2_FILL8
XSTDFILL106_680 VDD VSS sg13g2_FILL8
XSTDFILL106_688 VDD VSS sg13g2_FILL8
XSTDFILL106_696 VDD VSS sg13g2_FILL8
XSTDFILL106_704 VDD VSS sg13g2_FILL8
XSTDFILL106_712 VDD VSS sg13g2_FILL8
XSTDFILL106_720 VDD VSS sg13g2_FILL8
XSTDFILL106_728 VDD VSS sg13g2_FILL8
XSTDFILL106_736 VDD VSS sg13g2_FILL8
XSTDFILL106_744 VDD VSS sg13g2_FILL8
XSTDFILL106_752 VDD VSS sg13g2_FILL8
XSTDFILL106_760 VDD VSS sg13g2_FILL8
XSTDFILL106_768 VDD VSS sg13g2_FILL8
XSTDFILL106_776 VDD VSS sg13g2_FILL8
XSTDFILL106_784 VDD VSS sg13g2_FILL8
XSTDFILL106_792 VDD VSS sg13g2_FILL8
XSTDFILL106_800 VDD VSS sg13g2_FILL8
XSTDFILL106_808 VDD VSS sg13g2_FILL8
XSTDFILL106_816 VDD VSS sg13g2_FILL8
XSTDFILL106_824 VDD VSS sg13g2_FILL8
XSTDFILL106_832 VDD VSS sg13g2_FILL8
XSTDFILL106_840 VDD VSS sg13g2_FILL8
XSTDFILL106_848 VDD VSS sg13g2_FILL8
XSTDFILL106_856 VDD VSS sg13g2_FILL8
XSTDFILL106_864 VDD VSS sg13g2_FILL8
XSTDFILL106_872 VDD VSS sg13g2_FILL8
XSTDFILL106_880 VDD VSS sg13g2_FILL8
XSTDFILL106_888 VDD VSS sg13g2_FILL8
XSTDFILL106_896 VDD VSS sg13g2_FILL8
XSTDFILL106_904 VDD VSS sg13g2_FILL8
XSTDFILL106_912 VDD VSS sg13g2_FILL8
XSTDFILL106_920 VDD VSS sg13g2_FILL8
XSTDFILL106_928 VDD VSS sg13g2_FILL8
XSTDFILL106_936 VDD VSS sg13g2_FILL8
XSTDFILL106_944 VDD VSS sg13g2_FILL8
XSTDFILL106_952 VDD VSS sg13g2_FILL8
XSTDFILL106_960 VDD VSS sg13g2_FILL8
XSTDFILL106_968 VDD VSS sg13g2_FILL8
XSTDFILL106_976 VDD VSS sg13g2_FILL8
XSTDFILL106_984 VDD VSS sg13g2_FILL8
XSTDFILL106_992 VDD VSS sg13g2_FILL8
XSTDFILL106_1000 VDD VSS sg13g2_FILL8
XSTDFILL106_1008 VDD VSS sg13g2_FILL8
XSTDFILL106_1016 VDD VSS sg13g2_FILL8
XSTDFILL106_1024 VDD VSS sg13g2_FILL8
XSTDFILL106_1032 VDD VSS sg13g2_FILL8
XSTDFILL106_1040 VDD VSS sg13g2_FILL8
XSTDFILL106_1048 VDD VSS sg13g2_FILL8
XSTDFILL106_1056 VDD VSS sg13g2_FILL8
XSTDFILL106_1064 VDD VSS sg13g2_FILL8
XSTDFILL106_1072 VDD VSS sg13g2_FILL8
XSTDFILL106_1080 VDD VSS sg13g2_FILL8
XSTDFILL106_1088 VDD VSS sg13g2_FILL8
XSTDFILL106_1096 VDD VSS sg13g2_FILL8
XSTDFILL106_1104 VDD VSS sg13g2_FILL8
XSTDFILL106_1112 VDD VSS sg13g2_FILL8
XSTDFILL106_1120 VDD VSS sg13g2_FILL8
XSTDFILL106_1128 VDD VSS sg13g2_FILL8
XSTDFILL106_1136 VDD VSS sg13g2_FILL8
XSTDFILL106_1144 VDD VSS sg13g2_FILL8
XSTDFILL106_1152 VDD VSS sg13g2_FILL8
XSTDFILL106_1160 VDD VSS sg13g2_FILL8
XSTDFILL106_1168 VDD VSS sg13g2_FILL8
XSTDFILL106_1176 VDD VSS sg13g2_FILL8
XSTDFILL106_1184 VDD VSS sg13g2_FILL8
XSTDFILL106_1192 VDD VSS sg13g2_FILL8
XSTDFILL106_1200 VDD VSS sg13g2_FILL8
XSTDFILL106_1208 VDD VSS sg13g2_FILL8
XSTDFILL106_1216 VDD VSS sg13g2_FILL8
XSTDFILL106_1224 VDD VSS sg13g2_FILL8
XSTDFILL106_1232 VDD VSS sg13g2_FILL8
XSTDFILL106_1240 VDD VSS sg13g2_FILL8
XSTDFILL106_1248 VDD VSS sg13g2_FILL8
XSTDFILL106_1256 VDD VSS sg13g2_FILL8
XSTDFILL106_1264 VDD VSS sg13g2_FILL8
XSTDFILL106_1272 VDD VSS sg13g2_FILL8
XSTDFILL106_1280 VDD VSS sg13g2_FILL8
XSTDFILL106_1288 VDD VSS sg13g2_FILL8
XSTDFILL106_1296 VDD VSS sg13g2_FILL8
XSTDFILL106_1304 VDD VSS sg13g2_FILL8
XSTDFILL106_1312 VDD VSS sg13g2_FILL8
XSTDFILL106_1320 VDD VSS sg13g2_FILL8
XSTDFILL106_1328 VDD VSS sg13g2_FILL8
XSTDFILL106_1336 VDD VSS sg13g2_FILL8
XSTDFILL106_1344 VDD VSS sg13g2_FILL8
XSTDFILL106_1352 VDD VSS sg13g2_FILL8
XSTDFILL106_1360 VDD VSS sg13g2_FILL8
XSTDFILL106_1368 VDD VSS sg13g2_FILL8
XSTDFILL106_1376 VDD VSS sg13g2_FILL8
XSTDFILL106_1384 VDD VSS sg13g2_FILL8
XSTDFILL106_1392 VDD VSS sg13g2_FILL8
XSTDFILL106_1400 VDD VSS sg13g2_FILL8
XSTDFILL106_1408 VDD VSS sg13g2_FILL8
XSTDFILL106_1416 VDD VSS sg13g2_FILL8
XSTDFILL106_1424 VDD VSS sg13g2_FILL8
XSTDFILL106_1432 VDD VSS sg13g2_FILL8
XSTDFILL106_1440 VDD VSS sg13g2_FILL8
XSTDFILL106_1448 VDD VSS sg13g2_FILL8
XSTDFILL106_1456 VDD VSS sg13g2_FILL8
XSTDFILL106_1464 VDD VSS sg13g2_FILL8
XSTDFILL106_1472 VDD VSS sg13g2_FILL8
XSTDFILL106_1480 VDD VSS sg13g2_FILL8
XSTDFILL106_1488 VDD VSS sg13g2_FILL8
XSTDFILL106_1496 VDD VSS sg13g2_FILL8
XSTDFILL106_1504 VDD VSS sg13g2_FILL8
XSTDFILL106_1512 VDD VSS sg13g2_FILL8
XSTDFILL106_1520 VDD VSS sg13g2_FILL8
XSTDFILL106_1528 VDD VSS sg13g2_FILL2
XSTDFILL106_1530 VDD VSS sg13g2_FILL1
XSTDFILL107_0 VDD VSS sg13g2_FILL8
XSTDFILL107_8 VDD VSS sg13g2_FILL8
XSTDFILL107_16 VDD VSS sg13g2_FILL8
XSTDFILL107_24 VDD VSS sg13g2_FILL8
XSTDFILL107_32 VDD VSS sg13g2_FILL8
XSTDFILL107_40 VDD VSS sg13g2_FILL8
XSTDFILL107_48 VDD VSS sg13g2_FILL8
XSTDFILL107_56 VDD VSS sg13g2_FILL8
XSTDFILL107_64 VDD VSS sg13g2_FILL8
XSTDFILL107_72 VDD VSS sg13g2_FILL8
XSTDFILL107_80 VDD VSS sg13g2_FILL8
XSTDFILL107_88 VDD VSS sg13g2_FILL8
XSTDFILL107_96 VDD VSS sg13g2_FILL8
XSTDFILL107_104 VDD VSS sg13g2_FILL8
XSTDFILL107_112 VDD VSS sg13g2_FILL8
XSTDFILL107_120 VDD VSS sg13g2_FILL8
XSTDFILL107_128 VDD VSS sg13g2_FILL8
XSTDFILL107_136 VDD VSS sg13g2_FILL8
XSTDFILL107_144 VDD VSS sg13g2_FILL8
XSTDFILL107_152 VDD VSS sg13g2_FILL8
XSTDFILL107_160 VDD VSS sg13g2_FILL8
XSTDFILL107_168 VDD VSS sg13g2_FILL8
XSTDFILL107_176 VDD VSS sg13g2_FILL8
XSTDFILL107_184 VDD VSS sg13g2_FILL8
XSTDFILL107_192 VDD VSS sg13g2_FILL8
XSTDFILL107_200 VDD VSS sg13g2_FILL8
XSTDFILL107_208 VDD VSS sg13g2_FILL8
XSTDFILL107_216 VDD VSS sg13g2_FILL8
XSTDFILL107_224 VDD VSS sg13g2_FILL8
XSTDFILL107_232 VDD VSS sg13g2_FILL8
XSTDFILL107_240 VDD VSS sg13g2_FILL8
XSTDFILL107_248 VDD VSS sg13g2_FILL8
XSTDFILL107_256 VDD VSS sg13g2_FILL8
XSTDFILL107_264 VDD VSS sg13g2_FILL8
XSTDFILL107_272 VDD VSS sg13g2_FILL8
XSTDFILL107_280 VDD VSS sg13g2_FILL8
XSTDFILL107_288 VDD VSS sg13g2_FILL8
XSTDFILL107_296 VDD VSS sg13g2_FILL8
XSTDFILL107_304 VDD VSS sg13g2_FILL8
XSTDFILL107_312 VDD VSS sg13g2_FILL8
XSTDFILL107_320 VDD VSS sg13g2_FILL8
XSTDFILL107_328 VDD VSS sg13g2_FILL8
XSTDFILL107_336 VDD VSS sg13g2_FILL8
XSTDFILL107_344 VDD VSS sg13g2_FILL8
XSTDFILL107_352 VDD VSS sg13g2_FILL8
XSTDFILL107_360 VDD VSS sg13g2_FILL8
XSTDFILL107_368 VDD VSS sg13g2_FILL8
XSTDFILL107_376 VDD VSS sg13g2_FILL8
XSTDFILL107_384 VDD VSS sg13g2_FILL8
XSTDFILL107_392 VDD VSS sg13g2_FILL8
XSTDFILL107_400 VDD VSS sg13g2_FILL8
XSTDFILL107_408 VDD VSS sg13g2_FILL8
XSTDFILL107_416 VDD VSS sg13g2_FILL8
XSTDFILL107_424 VDD VSS sg13g2_FILL8
XSTDFILL107_432 VDD VSS sg13g2_FILL8
XSTDFILL107_440 VDD VSS sg13g2_FILL8
XSTDFILL107_448 VDD VSS sg13g2_FILL8
XSTDFILL107_456 VDD VSS sg13g2_FILL8
XSTDFILL107_464 VDD VSS sg13g2_FILL8
XSTDFILL107_472 VDD VSS sg13g2_FILL8
XSTDFILL107_480 VDD VSS sg13g2_FILL8
XSTDFILL107_488 VDD VSS sg13g2_FILL8
XSTDFILL107_496 VDD VSS sg13g2_FILL8
XSTDFILL107_504 VDD VSS sg13g2_FILL8
XSTDFILL107_512 VDD VSS sg13g2_FILL8
XSTDFILL107_520 VDD VSS sg13g2_FILL8
XSTDFILL107_528 VDD VSS sg13g2_FILL8
XSTDFILL107_536 VDD VSS sg13g2_FILL8
XSTDFILL107_544 VDD VSS sg13g2_FILL8
XSTDFILL107_552 VDD VSS sg13g2_FILL8
XSTDFILL107_560 VDD VSS sg13g2_FILL8
XSTDFILL107_568 VDD VSS sg13g2_FILL8
XSTDFILL107_576 VDD VSS sg13g2_FILL8
XSTDFILL107_584 VDD VSS sg13g2_FILL8
XSTDFILL107_592 VDD VSS sg13g2_FILL8
XSTDFILL107_600 VDD VSS sg13g2_FILL8
XSTDFILL107_608 VDD VSS sg13g2_FILL8
XSTDFILL107_616 VDD VSS sg13g2_FILL8
XSTDFILL107_624 VDD VSS sg13g2_FILL8
XSTDFILL107_632 VDD VSS sg13g2_FILL8
XSTDFILL107_640 VDD VSS sg13g2_FILL8
XSTDFILL107_648 VDD VSS sg13g2_FILL8
XSTDFILL107_656 VDD VSS sg13g2_FILL8
XSTDFILL107_664 VDD VSS sg13g2_FILL8
XSTDFILL107_672 VDD VSS sg13g2_FILL8
XSTDFILL107_680 VDD VSS sg13g2_FILL8
XSTDFILL107_688 VDD VSS sg13g2_FILL8
XSTDFILL107_696 VDD VSS sg13g2_FILL8
XSTDFILL107_704 VDD VSS sg13g2_FILL8
XSTDFILL107_712 VDD VSS sg13g2_FILL8
XSTDFILL107_720 VDD VSS sg13g2_FILL8
XSTDFILL107_728 VDD VSS sg13g2_FILL8
XSTDFILL107_736 VDD VSS sg13g2_FILL8
XSTDFILL107_744 VDD VSS sg13g2_FILL8
XSTDFILL107_752 VDD VSS sg13g2_FILL8
XSTDFILL107_760 VDD VSS sg13g2_FILL8
XSTDFILL107_768 VDD VSS sg13g2_FILL8
XSTDFILL107_776 VDD VSS sg13g2_FILL8
XSTDFILL107_784 VDD VSS sg13g2_FILL8
XSTDFILL107_792 VDD VSS sg13g2_FILL8
XSTDFILL107_800 VDD VSS sg13g2_FILL8
XSTDFILL107_808 VDD VSS sg13g2_FILL8
XSTDFILL107_816 VDD VSS sg13g2_FILL8
XSTDFILL107_824 VDD VSS sg13g2_FILL8
XSTDFILL107_832 VDD VSS sg13g2_FILL8
XSTDFILL107_840 VDD VSS sg13g2_FILL8
XSTDFILL107_848 VDD VSS sg13g2_FILL8
XSTDFILL107_856 VDD VSS sg13g2_FILL8
XSTDFILL107_864 VDD VSS sg13g2_FILL8
XSTDFILL107_872 VDD VSS sg13g2_FILL8
XSTDFILL107_880 VDD VSS sg13g2_FILL8
XSTDFILL107_888 VDD VSS sg13g2_FILL8
XSTDFILL107_896 VDD VSS sg13g2_FILL8
XSTDFILL107_904 VDD VSS sg13g2_FILL8
XSTDFILL107_912 VDD VSS sg13g2_FILL8
XSTDFILL107_920 VDD VSS sg13g2_FILL8
XSTDFILL107_928 VDD VSS sg13g2_FILL8
XSTDFILL107_936 VDD VSS sg13g2_FILL8
XSTDFILL107_944 VDD VSS sg13g2_FILL8
XSTDFILL107_952 VDD VSS sg13g2_FILL8
XSTDFILL107_960 VDD VSS sg13g2_FILL8
XSTDFILL107_968 VDD VSS sg13g2_FILL8
XSTDFILL107_976 VDD VSS sg13g2_FILL8
XSTDFILL107_984 VDD VSS sg13g2_FILL8
XSTDFILL107_992 VDD VSS sg13g2_FILL8
XSTDFILL107_1000 VDD VSS sg13g2_FILL8
XSTDFILL107_1008 VDD VSS sg13g2_FILL8
XSTDFILL107_1016 VDD VSS sg13g2_FILL8
XSTDFILL107_1024 VDD VSS sg13g2_FILL8
XSTDFILL107_1032 VDD VSS sg13g2_FILL8
XSTDFILL107_1040 VDD VSS sg13g2_FILL8
XSTDFILL107_1048 VDD VSS sg13g2_FILL8
XSTDFILL107_1056 VDD VSS sg13g2_FILL8
XSTDFILL107_1064 VDD VSS sg13g2_FILL8
XSTDFILL107_1072 VDD VSS sg13g2_FILL8
XSTDFILL107_1080 VDD VSS sg13g2_FILL8
XSTDFILL107_1088 VDD VSS sg13g2_FILL8
XSTDFILL107_1096 VDD VSS sg13g2_FILL8
XSTDFILL107_1104 VDD VSS sg13g2_FILL8
XSTDFILL107_1112 VDD VSS sg13g2_FILL8
XSTDFILL107_1120 VDD VSS sg13g2_FILL8
XSTDFILL107_1128 VDD VSS sg13g2_FILL8
XSTDFILL107_1136 VDD VSS sg13g2_FILL8
XSTDFILL107_1144 VDD VSS sg13g2_FILL8
XSTDFILL107_1152 VDD VSS sg13g2_FILL8
XSTDFILL107_1160 VDD VSS sg13g2_FILL8
XSTDFILL107_1168 VDD VSS sg13g2_FILL8
XSTDFILL107_1176 VDD VSS sg13g2_FILL8
XSTDFILL107_1184 VDD VSS sg13g2_FILL8
XSTDFILL107_1192 VDD VSS sg13g2_FILL8
XSTDFILL107_1200 VDD VSS sg13g2_FILL8
XSTDFILL107_1208 VDD VSS sg13g2_FILL8
XSTDFILL107_1216 VDD VSS sg13g2_FILL8
XSTDFILL107_1224 VDD VSS sg13g2_FILL8
XSTDFILL107_1232 VDD VSS sg13g2_FILL8
XSTDFILL107_1240 VDD VSS sg13g2_FILL8
XSTDFILL107_1248 VDD VSS sg13g2_FILL8
XSTDFILL107_1256 VDD VSS sg13g2_FILL8
XSTDFILL107_1264 VDD VSS sg13g2_FILL8
XSTDFILL107_1272 VDD VSS sg13g2_FILL8
XSTDFILL107_1280 VDD VSS sg13g2_FILL8
XSTDFILL107_1288 VDD VSS sg13g2_FILL8
XSTDFILL107_1296 VDD VSS sg13g2_FILL8
XSTDFILL107_1304 VDD VSS sg13g2_FILL8
XSTDFILL107_1312 VDD VSS sg13g2_FILL8
XSTDFILL107_1320 VDD VSS sg13g2_FILL8
XSTDFILL107_1328 VDD VSS sg13g2_FILL8
XSTDFILL107_1336 VDD VSS sg13g2_FILL8
XSTDFILL107_1344 VDD VSS sg13g2_FILL8
XSTDFILL107_1352 VDD VSS sg13g2_FILL8
XSTDFILL107_1360 VDD VSS sg13g2_FILL8
XSTDFILL107_1368 VDD VSS sg13g2_FILL8
XSTDFILL107_1376 VDD VSS sg13g2_FILL8
XSTDFILL107_1384 VDD VSS sg13g2_FILL8
XSTDFILL107_1392 VDD VSS sg13g2_FILL8
XSTDFILL107_1400 VDD VSS sg13g2_FILL8
XSTDFILL107_1408 VDD VSS sg13g2_FILL8
XSTDFILL107_1416 VDD VSS sg13g2_FILL8
XSTDFILL107_1424 VDD VSS sg13g2_FILL8
XSTDFILL107_1432 VDD VSS sg13g2_FILL8
XSTDFILL107_1440 VDD VSS sg13g2_FILL8
XSTDFILL107_1448 VDD VSS sg13g2_FILL8
XSTDFILL107_1456 VDD VSS sg13g2_FILL8
XSTDFILL107_1464 VDD VSS sg13g2_FILL8
XSTDFILL107_1472 VDD VSS sg13g2_FILL8
XSTDFILL107_1480 VDD VSS sg13g2_FILL8
XSTDFILL107_1488 VDD VSS sg13g2_FILL8
XSTDFILL107_1496 VDD VSS sg13g2_FILL8
XSTDFILL107_1504 VDD VSS sg13g2_FILL8
XSTDFILL107_1512 VDD VSS sg13g2_FILL8
XSTDFILL107_1520 VDD VSS sg13g2_FILL8
XSTDFILL107_1528 VDD VSS sg13g2_FILL2
XSTDFILL107_1530 VDD VSS sg13g2_FILL1
XSTDFILL108_0 VDD VSS sg13g2_FILL8
XSTDFILL108_8 VDD VSS sg13g2_FILL8
XSTDFILL108_16 VDD VSS sg13g2_FILL8
XSTDFILL108_24 VDD VSS sg13g2_FILL8
XSTDFILL108_32 VDD VSS sg13g2_FILL8
XSTDFILL108_40 VDD VSS sg13g2_FILL8
XSTDFILL108_48 VDD VSS sg13g2_FILL8
XSTDFILL108_56 VDD VSS sg13g2_FILL8
XSTDFILL108_64 VDD VSS sg13g2_FILL8
XSTDFILL108_72 VDD VSS sg13g2_FILL8
XSTDFILL108_80 VDD VSS sg13g2_FILL8
XSTDFILL108_88 VDD VSS sg13g2_FILL8
XSTDFILL108_96 VDD VSS sg13g2_FILL8
XSTDFILL108_104 VDD VSS sg13g2_FILL8
XSTDFILL108_112 VDD VSS sg13g2_FILL8
XSTDFILL108_120 VDD VSS sg13g2_FILL8
XSTDFILL108_128 VDD VSS sg13g2_FILL8
XSTDFILL108_136 VDD VSS sg13g2_FILL8
XSTDFILL108_144 VDD VSS sg13g2_FILL8
XSTDFILL108_152 VDD VSS sg13g2_FILL8
XSTDFILL108_160 VDD VSS sg13g2_FILL8
XSTDFILL108_168 VDD VSS sg13g2_FILL8
XSTDFILL108_176 VDD VSS sg13g2_FILL8
XSTDFILL108_184 VDD VSS sg13g2_FILL8
XSTDFILL108_192 VDD VSS sg13g2_FILL8
XSTDFILL108_200 VDD VSS sg13g2_FILL8
XSTDFILL108_208 VDD VSS sg13g2_FILL8
XSTDFILL108_216 VDD VSS sg13g2_FILL8
XSTDFILL108_224 VDD VSS sg13g2_FILL8
XSTDFILL108_232 VDD VSS sg13g2_FILL8
XSTDFILL108_240 VDD VSS sg13g2_FILL8
XSTDFILL108_248 VDD VSS sg13g2_FILL8
XSTDFILL108_256 VDD VSS sg13g2_FILL8
XSTDFILL108_264 VDD VSS sg13g2_FILL8
XSTDFILL108_272 VDD VSS sg13g2_FILL8
XSTDFILL108_280 VDD VSS sg13g2_FILL8
XSTDFILL108_288 VDD VSS sg13g2_FILL8
XSTDFILL108_296 VDD VSS sg13g2_FILL8
XSTDFILL108_304 VDD VSS sg13g2_FILL8
XSTDFILL108_312 VDD VSS sg13g2_FILL8
XSTDFILL108_320 VDD VSS sg13g2_FILL8
XSTDFILL108_328 VDD VSS sg13g2_FILL8
XSTDFILL108_336 VDD VSS sg13g2_FILL8
XSTDFILL108_344 VDD VSS sg13g2_FILL8
XSTDFILL108_352 VDD VSS sg13g2_FILL8
XSTDFILL108_360 VDD VSS sg13g2_FILL8
XSTDFILL108_368 VDD VSS sg13g2_FILL8
XSTDFILL108_376 VDD VSS sg13g2_FILL8
XSTDFILL108_384 VDD VSS sg13g2_FILL8
XSTDFILL108_392 VDD VSS sg13g2_FILL8
XSTDFILL108_400 VDD VSS sg13g2_FILL8
XSTDFILL108_408 VDD VSS sg13g2_FILL8
XSTDFILL108_416 VDD VSS sg13g2_FILL8
XSTDFILL108_424 VDD VSS sg13g2_FILL8
XSTDFILL108_432 VDD VSS sg13g2_FILL8
XSTDFILL108_440 VDD VSS sg13g2_FILL8
XSTDFILL108_448 VDD VSS sg13g2_FILL8
XSTDFILL108_456 VDD VSS sg13g2_FILL8
XSTDFILL108_464 VDD VSS sg13g2_FILL8
XSTDFILL108_472 VDD VSS sg13g2_FILL8
XSTDFILL108_480 VDD VSS sg13g2_FILL8
XSTDFILL108_488 VDD VSS sg13g2_FILL8
XSTDFILL108_496 VDD VSS sg13g2_FILL8
XSTDFILL108_504 VDD VSS sg13g2_FILL8
XSTDFILL108_512 VDD VSS sg13g2_FILL8
XSTDFILL108_520 VDD VSS sg13g2_FILL8
XSTDFILL108_528 VDD VSS sg13g2_FILL8
XSTDFILL108_536 VDD VSS sg13g2_FILL8
XSTDFILL108_544 VDD VSS sg13g2_FILL8
XSTDFILL108_552 VDD VSS sg13g2_FILL8
XSTDFILL108_560 VDD VSS sg13g2_FILL8
XSTDFILL108_568 VDD VSS sg13g2_FILL8
XSTDFILL108_576 VDD VSS sg13g2_FILL8
XSTDFILL108_584 VDD VSS sg13g2_FILL8
XSTDFILL108_592 VDD VSS sg13g2_FILL8
XSTDFILL108_600 VDD VSS sg13g2_FILL8
XSTDFILL108_608 VDD VSS sg13g2_FILL8
XSTDFILL108_616 VDD VSS sg13g2_FILL8
XSTDFILL108_624 VDD VSS sg13g2_FILL8
XSTDFILL108_632 VDD VSS sg13g2_FILL8
XSTDFILL108_640 VDD VSS sg13g2_FILL8
XSTDFILL108_648 VDD VSS sg13g2_FILL8
XSTDFILL108_656 VDD VSS sg13g2_FILL8
XSTDFILL108_664 VDD VSS sg13g2_FILL8
XSTDFILL108_672 VDD VSS sg13g2_FILL8
XSTDFILL108_680 VDD VSS sg13g2_FILL8
XSTDFILL108_688 VDD VSS sg13g2_FILL8
XSTDFILL108_696 VDD VSS sg13g2_FILL8
XSTDFILL108_704 VDD VSS sg13g2_FILL8
XSTDFILL108_712 VDD VSS sg13g2_FILL8
XSTDFILL108_720 VDD VSS sg13g2_FILL8
XSTDFILL108_728 VDD VSS sg13g2_FILL8
XSTDFILL108_736 VDD VSS sg13g2_FILL8
XSTDFILL108_744 VDD VSS sg13g2_FILL8
XSTDFILL108_752 VDD VSS sg13g2_FILL8
XSTDFILL108_760 VDD VSS sg13g2_FILL8
XSTDFILL108_768 VDD VSS sg13g2_FILL8
XSTDFILL108_776 VDD VSS sg13g2_FILL8
XSTDFILL108_784 VDD VSS sg13g2_FILL8
XSTDFILL108_792 VDD VSS sg13g2_FILL8
XSTDFILL108_800 VDD VSS sg13g2_FILL8
XSTDFILL108_808 VDD VSS sg13g2_FILL8
XSTDFILL108_816 VDD VSS sg13g2_FILL8
XSTDFILL108_824 VDD VSS sg13g2_FILL8
XSTDFILL108_832 VDD VSS sg13g2_FILL8
XSTDFILL108_840 VDD VSS sg13g2_FILL8
XSTDFILL108_848 VDD VSS sg13g2_FILL8
XSTDFILL108_856 VDD VSS sg13g2_FILL8
XSTDFILL108_864 VDD VSS sg13g2_FILL8
XSTDFILL108_872 VDD VSS sg13g2_FILL8
XSTDFILL108_880 VDD VSS sg13g2_FILL8
XSTDFILL108_888 VDD VSS sg13g2_FILL8
XSTDFILL108_896 VDD VSS sg13g2_FILL8
XSTDFILL108_904 VDD VSS sg13g2_FILL8
XSTDFILL108_912 VDD VSS sg13g2_FILL8
XSTDFILL108_920 VDD VSS sg13g2_FILL8
XSTDFILL108_928 VDD VSS sg13g2_FILL8
XSTDFILL108_936 VDD VSS sg13g2_FILL8
XSTDFILL108_944 VDD VSS sg13g2_FILL8
XSTDFILL108_952 VDD VSS sg13g2_FILL8
XSTDFILL108_960 VDD VSS sg13g2_FILL8
XSTDFILL108_968 VDD VSS sg13g2_FILL8
XSTDFILL108_976 VDD VSS sg13g2_FILL8
XSTDFILL108_984 VDD VSS sg13g2_FILL8
XSTDFILL108_992 VDD VSS sg13g2_FILL8
XSTDFILL108_1000 VDD VSS sg13g2_FILL8
XSTDFILL108_1008 VDD VSS sg13g2_FILL8
XSTDFILL108_1016 VDD VSS sg13g2_FILL8
XSTDFILL108_1024 VDD VSS sg13g2_FILL8
XSTDFILL108_1032 VDD VSS sg13g2_FILL8
XSTDFILL108_1040 VDD VSS sg13g2_FILL8
XSTDFILL108_1048 VDD VSS sg13g2_FILL8
XSTDFILL108_1056 VDD VSS sg13g2_FILL8
XSTDFILL108_1064 VDD VSS sg13g2_FILL8
XSTDFILL108_1072 VDD VSS sg13g2_FILL8
XSTDFILL108_1080 VDD VSS sg13g2_FILL8
XSTDFILL108_1088 VDD VSS sg13g2_FILL8
XSTDFILL108_1096 VDD VSS sg13g2_FILL8
XSTDFILL108_1104 VDD VSS sg13g2_FILL8
XSTDFILL108_1112 VDD VSS sg13g2_FILL8
XSTDFILL108_1120 VDD VSS sg13g2_FILL8
XSTDFILL108_1128 VDD VSS sg13g2_FILL8
XSTDFILL108_1136 VDD VSS sg13g2_FILL8
XSTDFILL108_1144 VDD VSS sg13g2_FILL8
XSTDFILL108_1152 VDD VSS sg13g2_FILL8
XSTDFILL108_1160 VDD VSS sg13g2_FILL8
XSTDFILL108_1168 VDD VSS sg13g2_FILL8
XSTDFILL108_1176 VDD VSS sg13g2_FILL8
XSTDFILL108_1184 VDD VSS sg13g2_FILL8
XSTDFILL108_1192 VDD VSS sg13g2_FILL8
XSTDFILL108_1200 VDD VSS sg13g2_FILL8
XSTDFILL108_1208 VDD VSS sg13g2_FILL8
XSTDFILL108_1216 VDD VSS sg13g2_FILL8
XSTDFILL108_1224 VDD VSS sg13g2_FILL8
XSTDFILL108_1232 VDD VSS sg13g2_FILL8
XSTDFILL108_1240 VDD VSS sg13g2_FILL8
XSTDFILL108_1248 VDD VSS sg13g2_FILL8
XSTDFILL108_1256 VDD VSS sg13g2_FILL8
XSTDFILL108_1264 VDD VSS sg13g2_FILL8
XSTDFILL108_1272 VDD VSS sg13g2_FILL8
XSTDFILL108_1280 VDD VSS sg13g2_FILL8
XSTDFILL108_1288 VDD VSS sg13g2_FILL8
XSTDFILL108_1296 VDD VSS sg13g2_FILL8
XSTDFILL108_1304 VDD VSS sg13g2_FILL8
XSTDFILL108_1312 VDD VSS sg13g2_FILL8
XSTDFILL108_1320 VDD VSS sg13g2_FILL8
XSTDFILL108_1328 VDD VSS sg13g2_FILL8
XSTDFILL108_1336 VDD VSS sg13g2_FILL8
XSTDFILL108_1344 VDD VSS sg13g2_FILL8
XSTDFILL108_1352 VDD VSS sg13g2_FILL8
XSTDFILL108_1360 VDD VSS sg13g2_FILL8
XSTDFILL108_1368 VDD VSS sg13g2_FILL8
XSTDFILL108_1376 VDD VSS sg13g2_FILL8
XSTDFILL108_1384 VDD VSS sg13g2_FILL8
XSTDFILL108_1392 VDD VSS sg13g2_FILL8
XSTDFILL108_1400 VDD VSS sg13g2_FILL8
XSTDFILL108_1408 VDD VSS sg13g2_FILL8
XSTDFILL108_1416 VDD VSS sg13g2_FILL8
XSTDFILL108_1424 VDD VSS sg13g2_FILL8
XSTDFILL108_1432 VDD VSS sg13g2_FILL8
XSTDFILL108_1440 VDD VSS sg13g2_FILL8
XSTDFILL108_1448 VDD VSS sg13g2_FILL8
XSTDFILL108_1456 VDD VSS sg13g2_FILL8
XSTDFILL108_1464 VDD VSS sg13g2_FILL8
XSTDFILL108_1472 VDD VSS sg13g2_FILL8
XSTDFILL108_1480 VDD VSS sg13g2_FILL8
XSTDFILL108_1488 VDD VSS sg13g2_FILL8
XSTDFILL108_1496 VDD VSS sg13g2_FILL8
XSTDFILL108_1504 VDD VSS sg13g2_FILL8
XSTDFILL108_1512 VDD VSS sg13g2_FILL8
XSTDFILL108_1520 VDD VSS sg13g2_FILL8
XSTDFILL108_1528 VDD VSS sg13g2_FILL2
XSTDFILL108_1530 VDD VSS sg13g2_FILL1
XSTDFILL109_0 VDD VSS sg13g2_FILL8
XSTDFILL109_8 VDD VSS sg13g2_FILL8
XSTDFILL109_16 VDD VSS sg13g2_FILL8
XSTDFILL109_24 VDD VSS sg13g2_FILL8
XSTDFILL109_32 VDD VSS sg13g2_FILL8
XSTDFILL109_40 VDD VSS sg13g2_FILL8
XSTDFILL109_48 VDD VSS sg13g2_FILL8
XSTDFILL109_56 VDD VSS sg13g2_FILL8
XSTDFILL109_64 VDD VSS sg13g2_FILL8
XSTDFILL109_72 VDD VSS sg13g2_FILL8
XSTDFILL109_80 VDD VSS sg13g2_FILL8
XSTDFILL109_88 VDD VSS sg13g2_FILL8
XSTDFILL109_96 VDD VSS sg13g2_FILL8
XSTDFILL109_104 VDD VSS sg13g2_FILL8
XSTDFILL109_112 VDD VSS sg13g2_FILL8
XSTDFILL109_120 VDD VSS sg13g2_FILL8
XSTDFILL109_128 VDD VSS sg13g2_FILL8
XSTDFILL109_136 VDD VSS sg13g2_FILL8
XSTDFILL109_144 VDD VSS sg13g2_FILL8
XSTDFILL109_152 VDD VSS sg13g2_FILL8
XSTDFILL109_160 VDD VSS sg13g2_FILL8
XSTDFILL109_168 VDD VSS sg13g2_FILL8
XSTDFILL109_176 VDD VSS sg13g2_FILL8
XSTDFILL109_184 VDD VSS sg13g2_FILL8
XSTDFILL109_192 VDD VSS sg13g2_FILL8
XSTDFILL109_200 VDD VSS sg13g2_FILL8
XSTDFILL109_208 VDD VSS sg13g2_FILL8
XSTDFILL109_216 VDD VSS sg13g2_FILL8
XSTDFILL109_224 VDD VSS sg13g2_FILL8
XSTDFILL109_232 VDD VSS sg13g2_FILL8
XSTDFILL109_240 VDD VSS sg13g2_FILL8
XSTDFILL109_248 VDD VSS sg13g2_FILL8
XSTDFILL109_256 VDD VSS sg13g2_FILL8
XSTDFILL109_264 VDD VSS sg13g2_FILL8
XSTDFILL109_272 VDD VSS sg13g2_FILL8
XSTDFILL109_280 VDD VSS sg13g2_FILL8
XSTDFILL109_288 VDD VSS sg13g2_FILL8
XSTDFILL109_296 VDD VSS sg13g2_FILL8
XSTDFILL109_304 VDD VSS sg13g2_FILL8
XSTDFILL109_312 VDD VSS sg13g2_FILL8
XSTDFILL109_320 VDD VSS sg13g2_FILL8
XSTDFILL109_328 VDD VSS sg13g2_FILL8
XSTDFILL109_336 VDD VSS sg13g2_FILL8
XSTDFILL109_344 VDD VSS sg13g2_FILL8
XSTDFILL109_352 VDD VSS sg13g2_FILL8
XSTDFILL109_360 VDD VSS sg13g2_FILL8
XSTDFILL109_368 VDD VSS sg13g2_FILL8
XSTDFILL109_376 VDD VSS sg13g2_FILL8
XSTDFILL109_384 VDD VSS sg13g2_FILL8
XSTDFILL109_392 VDD VSS sg13g2_FILL8
XSTDFILL109_400 VDD VSS sg13g2_FILL8
XSTDFILL109_408 VDD VSS sg13g2_FILL8
XSTDFILL109_416 VDD VSS sg13g2_FILL8
XSTDFILL109_424 VDD VSS sg13g2_FILL8
XSTDFILL109_432 VDD VSS sg13g2_FILL8
XSTDFILL109_440 VDD VSS sg13g2_FILL8
XSTDFILL109_448 VDD VSS sg13g2_FILL8
XSTDFILL109_456 VDD VSS sg13g2_FILL8
XSTDFILL109_464 VDD VSS sg13g2_FILL8
XSTDFILL109_472 VDD VSS sg13g2_FILL8
XSTDFILL109_480 VDD VSS sg13g2_FILL8
XSTDFILL109_488 VDD VSS sg13g2_FILL8
XSTDFILL109_496 VDD VSS sg13g2_FILL8
XSTDFILL109_504 VDD VSS sg13g2_FILL8
XSTDFILL109_512 VDD VSS sg13g2_FILL8
XSTDFILL109_520 VDD VSS sg13g2_FILL8
XSTDFILL109_528 VDD VSS sg13g2_FILL8
XSTDFILL109_536 VDD VSS sg13g2_FILL8
XSTDFILL109_544 VDD VSS sg13g2_FILL8
XSTDFILL109_552 VDD VSS sg13g2_FILL8
XSTDFILL109_560 VDD VSS sg13g2_FILL8
XSTDFILL109_568 VDD VSS sg13g2_FILL8
XSTDFILL109_576 VDD VSS sg13g2_FILL8
XSTDFILL109_584 VDD VSS sg13g2_FILL8
XSTDFILL109_592 VDD VSS sg13g2_FILL8
XSTDFILL109_600 VDD VSS sg13g2_FILL8
XSTDFILL109_608 VDD VSS sg13g2_FILL8
XSTDFILL109_616 VDD VSS sg13g2_FILL8
XSTDFILL109_624 VDD VSS sg13g2_FILL8
XSTDFILL109_632 VDD VSS sg13g2_FILL8
XSTDFILL109_640 VDD VSS sg13g2_FILL8
XSTDFILL109_648 VDD VSS sg13g2_FILL8
XSTDFILL109_656 VDD VSS sg13g2_FILL8
XSTDFILL109_664 VDD VSS sg13g2_FILL8
XSTDFILL109_672 VDD VSS sg13g2_FILL8
XSTDFILL109_680 VDD VSS sg13g2_FILL8
XSTDFILL109_688 VDD VSS sg13g2_FILL8
XSTDFILL109_696 VDD VSS sg13g2_FILL8
XSTDFILL109_704 VDD VSS sg13g2_FILL8
XSTDFILL109_712 VDD VSS sg13g2_FILL8
XSTDFILL109_720 VDD VSS sg13g2_FILL8
XSTDFILL109_728 VDD VSS sg13g2_FILL8
XSTDFILL109_736 VDD VSS sg13g2_FILL8
XSTDFILL109_744 VDD VSS sg13g2_FILL8
XSTDFILL109_752 VDD VSS sg13g2_FILL8
XSTDFILL109_760 VDD VSS sg13g2_FILL8
XSTDFILL109_768 VDD VSS sg13g2_FILL8
XSTDFILL109_776 VDD VSS sg13g2_FILL8
XSTDFILL109_784 VDD VSS sg13g2_FILL8
XSTDFILL109_792 VDD VSS sg13g2_FILL8
XSTDFILL109_800 VDD VSS sg13g2_FILL8
XSTDFILL109_808 VDD VSS sg13g2_FILL8
XSTDFILL109_816 VDD VSS sg13g2_FILL8
XSTDFILL109_824 VDD VSS sg13g2_FILL8
XSTDFILL109_832 VDD VSS sg13g2_FILL8
XSTDFILL109_840 VDD VSS sg13g2_FILL8
XSTDFILL109_848 VDD VSS sg13g2_FILL8
XSTDFILL109_856 VDD VSS sg13g2_FILL8
XSTDFILL109_864 VDD VSS sg13g2_FILL8
XSTDFILL109_872 VDD VSS sg13g2_FILL8
XSTDFILL109_880 VDD VSS sg13g2_FILL8
XSTDFILL109_888 VDD VSS sg13g2_FILL8
XSTDFILL109_896 VDD VSS sg13g2_FILL8
XSTDFILL109_904 VDD VSS sg13g2_FILL8
XSTDFILL109_912 VDD VSS sg13g2_FILL8
XSTDFILL109_920 VDD VSS sg13g2_FILL8
XSTDFILL109_928 VDD VSS sg13g2_FILL8
XSTDFILL109_936 VDD VSS sg13g2_FILL8
XSTDFILL109_944 VDD VSS sg13g2_FILL8
XSTDFILL109_952 VDD VSS sg13g2_FILL8
XSTDFILL109_960 VDD VSS sg13g2_FILL8
XSTDFILL109_968 VDD VSS sg13g2_FILL8
XSTDFILL109_976 VDD VSS sg13g2_FILL8
XSTDFILL109_984 VDD VSS sg13g2_FILL8
XSTDFILL109_992 VDD VSS sg13g2_FILL8
XSTDFILL109_1000 VDD VSS sg13g2_FILL8
XSTDFILL109_1008 VDD VSS sg13g2_FILL8
XSTDFILL109_1016 VDD VSS sg13g2_FILL8
XSTDFILL109_1024 VDD VSS sg13g2_FILL8
XSTDFILL109_1032 VDD VSS sg13g2_FILL8
XSTDFILL109_1040 VDD VSS sg13g2_FILL8
XSTDFILL109_1048 VDD VSS sg13g2_FILL8
XSTDFILL109_1056 VDD VSS sg13g2_FILL8
XSTDFILL109_1064 VDD VSS sg13g2_FILL8
XSTDFILL109_1072 VDD VSS sg13g2_FILL8
XSTDFILL109_1080 VDD VSS sg13g2_FILL8
XSTDFILL109_1088 VDD VSS sg13g2_FILL8
XSTDFILL109_1096 VDD VSS sg13g2_FILL8
XSTDFILL109_1104 VDD VSS sg13g2_FILL8
XSTDFILL109_1112 VDD VSS sg13g2_FILL8
XSTDFILL109_1120 VDD VSS sg13g2_FILL8
XSTDFILL109_1128 VDD VSS sg13g2_FILL8
XSTDFILL109_1136 VDD VSS sg13g2_FILL8
XSTDFILL109_1144 VDD VSS sg13g2_FILL8
XSTDFILL109_1152 VDD VSS sg13g2_FILL8
XSTDFILL109_1160 VDD VSS sg13g2_FILL8
XSTDFILL109_1168 VDD VSS sg13g2_FILL8
XSTDFILL109_1176 VDD VSS sg13g2_FILL8
XSTDFILL109_1184 VDD VSS sg13g2_FILL8
XSTDFILL109_1192 VDD VSS sg13g2_FILL8
XSTDFILL109_1200 VDD VSS sg13g2_FILL8
XSTDFILL109_1208 VDD VSS sg13g2_FILL8
XSTDFILL109_1216 VDD VSS sg13g2_FILL8
XSTDFILL109_1224 VDD VSS sg13g2_FILL8
XSTDFILL109_1232 VDD VSS sg13g2_FILL8
XSTDFILL109_1240 VDD VSS sg13g2_FILL8
XSTDFILL109_1248 VDD VSS sg13g2_FILL8
XSTDFILL109_1256 VDD VSS sg13g2_FILL8
XSTDFILL109_1264 VDD VSS sg13g2_FILL8
XSTDFILL109_1272 VDD VSS sg13g2_FILL8
XSTDFILL109_1280 VDD VSS sg13g2_FILL8
XSTDFILL109_1288 VDD VSS sg13g2_FILL8
XSTDFILL109_1296 VDD VSS sg13g2_FILL8
XSTDFILL109_1304 VDD VSS sg13g2_FILL8
XSTDFILL109_1312 VDD VSS sg13g2_FILL8
XSTDFILL109_1320 VDD VSS sg13g2_FILL8
XSTDFILL109_1328 VDD VSS sg13g2_FILL8
XSTDFILL109_1336 VDD VSS sg13g2_FILL8
XSTDFILL109_1344 VDD VSS sg13g2_FILL8
XSTDFILL109_1352 VDD VSS sg13g2_FILL8
XSTDFILL109_1360 VDD VSS sg13g2_FILL8
XSTDFILL109_1368 VDD VSS sg13g2_FILL8
XSTDFILL109_1376 VDD VSS sg13g2_FILL8
XSTDFILL109_1384 VDD VSS sg13g2_FILL8
XSTDFILL109_1392 VDD VSS sg13g2_FILL8
XSTDFILL109_1400 VDD VSS sg13g2_FILL8
XSTDFILL109_1408 VDD VSS sg13g2_FILL8
XSTDFILL109_1416 VDD VSS sg13g2_FILL8
XSTDFILL109_1424 VDD VSS sg13g2_FILL8
XSTDFILL109_1432 VDD VSS sg13g2_FILL8
XSTDFILL109_1440 VDD VSS sg13g2_FILL8
XSTDFILL109_1448 VDD VSS sg13g2_FILL8
XSTDFILL109_1456 VDD VSS sg13g2_FILL8
XSTDFILL109_1464 VDD VSS sg13g2_FILL8
XSTDFILL109_1472 VDD VSS sg13g2_FILL8
XSTDFILL109_1480 VDD VSS sg13g2_FILL8
XSTDFILL109_1488 VDD VSS sg13g2_FILL8
XSTDFILL109_1496 VDD VSS sg13g2_FILL8
XSTDFILL109_1504 VDD VSS sg13g2_FILL8
XSTDFILL109_1512 VDD VSS sg13g2_FILL8
XSTDFILL109_1520 VDD VSS sg13g2_FILL8
XSTDFILL109_1528 VDD VSS sg13g2_FILL2
XSTDFILL109_1530 VDD VSS sg13g2_FILL1
XSTDFILL110_0 VDD VSS sg13g2_FILL8
XSTDFILL110_8 VDD VSS sg13g2_FILL8
XSTDFILL110_16 VDD VSS sg13g2_FILL8
XSTDFILL110_24 VDD VSS sg13g2_FILL8
XSTDFILL110_32 VDD VSS sg13g2_FILL8
XSTDFILL110_40 VDD VSS sg13g2_FILL8
XSTDFILL110_48 VDD VSS sg13g2_FILL8
XSTDFILL110_56 VDD VSS sg13g2_FILL8
XSTDFILL110_64 VDD VSS sg13g2_FILL8
XSTDFILL110_72 VDD VSS sg13g2_FILL8
XSTDFILL110_80 VDD VSS sg13g2_FILL8
XSTDFILL110_88 VDD VSS sg13g2_FILL8
XSTDFILL110_96 VDD VSS sg13g2_FILL8
XSTDFILL110_104 VDD VSS sg13g2_FILL8
XSTDFILL110_112 VDD VSS sg13g2_FILL8
XSTDFILL110_120 VDD VSS sg13g2_FILL8
XSTDFILL110_128 VDD VSS sg13g2_FILL8
XSTDFILL110_136 VDD VSS sg13g2_FILL8
XSTDFILL110_144 VDD VSS sg13g2_FILL8
XSTDFILL110_152 VDD VSS sg13g2_FILL8
XSTDFILL110_160 VDD VSS sg13g2_FILL8
XSTDFILL110_168 VDD VSS sg13g2_FILL8
XSTDFILL110_176 VDD VSS sg13g2_FILL8
XSTDFILL110_184 VDD VSS sg13g2_FILL8
XSTDFILL110_192 VDD VSS sg13g2_FILL8
XSTDFILL110_200 VDD VSS sg13g2_FILL8
XSTDFILL110_208 VDD VSS sg13g2_FILL8
XSTDFILL110_216 VDD VSS sg13g2_FILL8
XSTDFILL110_224 VDD VSS sg13g2_FILL8
XSTDFILL110_232 VDD VSS sg13g2_FILL8
XSTDFILL110_240 VDD VSS sg13g2_FILL8
XSTDFILL110_248 VDD VSS sg13g2_FILL8
XSTDFILL110_256 VDD VSS sg13g2_FILL8
XSTDFILL110_264 VDD VSS sg13g2_FILL8
XSTDFILL110_272 VDD VSS sg13g2_FILL8
XSTDFILL110_280 VDD VSS sg13g2_FILL8
XSTDFILL110_288 VDD VSS sg13g2_FILL8
XSTDFILL110_296 VDD VSS sg13g2_FILL8
XSTDFILL110_304 VDD VSS sg13g2_FILL8
XSTDFILL110_312 VDD VSS sg13g2_FILL8
XSTDFILL110_320 VDD VSS sg13g2_FILL8
XSTDFILL110_328 VDD VSS sg13g2_FILL8
XSTDFILL110_336 VDD VSS sg13g2_FILL8
XSTDFILL110_344 VDD VSS sg13g2_FILL8
XSTDFILL110_352 VDD VSS sg13g2_FILL8
XSTDFILL110_360 VDD VSS sg13g2_FILL8
XSTDFILL110_368 VDD VSS sg13g2_FILL8
XSTDFILL110_376 VDD VSS sg13g2_FILL8
XSTDFILL110_384 VDD VSS sg13g2_FILL8
XSTDFILL110_392 VDD VSS sg13g2_FILL8
XSTDFILL110_400 VDD VSS sg13g2_FILL8
XSTDFILL110_408 VDD VSS sg13g2_FILL8
XSTDFILL110_416 VDD VSS sg13g2_FILL8
XSTDFILL110_424 VDD VSS sg13g2_FILL8
XSTDFILL110_432 VDD VSS sg13g2_FILL8
XSTDFILL110_440 VDD VSS sg13g2_FILL8
XSTDFILL110_448 VDD VSS sg13g2_FILL8
XSTDFILL110_456 VDD VSS sg13g2_FILL8
XSTDFILL110_464 VDD VSS sg13g2_FILL8
XSTDFILL110_472 VDD VSS sg13g2_FILL8
XSTDFILL110_480 VDD VSS sg13g2_FILL8
XSTDFILL110_488 VDD VSS sg13g2_FILL8
XSTDFILL110_496 VDD VSS sg13g2_FILL8
XSTDFILL110_504 VDD VSS sg13g2_FILL8
XSTDFILL110_512 VDD VSS sg13g2_FILL8
XSTDFILL110_520 VDD VSS sg13g2_FILL8
XSTDFILL110_528 VDD VSS sg13g2_FILL8
XSTDFILL110_536 VDD VSS sg13g2_FILL8
XSTDFILL110_544 VDD VSS sg13g2_FILL8
XSTDFILL110_552 VDD VSS sg13g2_FILL8
XSTDFILL110_560 VDD VSS sg13g2_FILL8
XSTDFILL110_568 VDD VSS sg13g2_FILL8
XSTDFILL110_576 VDD VSS sg13g2_FILL8
XSTDFILL110_584 VDD VSS sg13g2_FILL8
XSTDFILL110_592 VDD VSS sg13g2_FILL8
XSTDFILL110_600 VDD VSS sg13g2_FILL8
XSTDFILL110_608 VDD VSS sg13g2_FILL8
XSTDFILL110_616 VDD VSS sg13g2_FILL8
XSTDFILL110_624 VDD VSS sg13g2_FILL8
XSTDFILL110_632 VDD VSS sg13g2_FILL8
XSTDFILL110_640 VDD VSS sg13g2_FILL8
XSTDFILL110_648 VDD VSS sg13g2_FILL8
XSTDFILL110_656 VDD VSS sg13g2_FILL8
XSTDFILL110_664 VDD VSS sg13g2_FILL8
XSTDFILL110_672 VDD VSS sg13g2_FILL8
XSTDFILL110_680 VDD VSS sg13g2_FILL8
XSTDFILL110_688 VDD VSS sg13g2_FILL8
XSTDFILL110_696 VDD VSS sg13g2_FILL8
XSTDFILL110_704 VDD VSS sg13g2_FILL8
XSTDFILL110_712 VDD VSS sg13g2_FILL8
XSTDFILL110_720 VDD VSS sg13g2_FILL8
XSTDFILL110_728 VDD VSS sg13g2_FILL8
XSTDFILL110_736 VDD VSS sg13g2_FILL8
XSTDFILL110_744 VDD VSS sg13g2_FILL8
XSTDFILL110_752 VDD VSS sg13g2_FILL8
XSTDFILL110_760 VDD VSS sg13g2_FILL8
XSTDFILL110_768 VDD VSS sg13g2_FILL8
XSTDFILL110_776 VDD VSS sg13g2_FILL8
XSTDFILL110_784 VDD VSS sg13g2_FILL8
XSTDFILL110_792 VDD VSS sg13g2_FILL8
XSTDFILL110_800 VDD VSS sg13g2_FILL8
XSTDFILL110_808 VDD VSS sg13g2_FILL8
XSTDFILL110_816 VDD VSS sg13g2_FILL8
XSTDFILL110_824 VDD VSS sg13g2_FILL8
XSTDFILL110_832 VDD VSS sg13g2_FILL8
XSTDFILL110_840 VDD VSS sg13g2_FILL8
XSTDFILL110_848 VDD VSS sg13g2_FILL8
XSTDFILL110_856 VDD VSS sg13g2_FILL8
XSTDFILL110_864 VDD VSS sg13g2_FILL8
XSTDFILL110_872 VDD VSS sg13g2_FILL8
XSTDFILL110_880 VDD VSS sg13g2_FILL8
XSTDFILL110_888 VDD VSS sg13g2_FILL8
XSTDFILL110_896 VDD VSS sg13g2_FILL8
XSTDFILL110_904 VDD VSS sg13g2_FILL8
XSTDFILL110_912 VDD VSS sg13g2_FILL8
XSTDFILL110_920 VDD VSS sg13g2_FILL8
XSTDFILL110_928 VDD VSS sg13g2_FILL8
XSTDFILL110_936 VDD VSS sg13g2_FILL8
XSTDFILL110_944 VDD VSS sg13g2_FILL8
XSTDFILL110_952 VDD VSS sg13g2_FILL8
XSTDFILL110_960 VDD VSS sg13g2_FILL8
XSTDFILL110_968 VDD VSS sg13g2_FILL8
XSTDFILL110_976 VDD VSS sg13g2_FILL8
XSTDFILL110_984 VDD VSS sg13g2_FILL8
XSTDFILL110_992 VDD VSS sg13g2_FILL8
XSTDFILL110_1000 VDD VSS sg13g2_FILL8
XSTDFILL110_1008 VDD VSS sg13g2_FILL8
XSTDFILL110_1016 VDD VSS sg13g2_FILL8
XSTDFILL110_1024 VDD VSS sg13g2_FILL8
XSTDFILL110_1032 VDD VSS sg13g2_FILL8
XSTDFILL110_1040 VDD VSS sg13g2_FILL8
XSTDFILL110_1048 VDD VSS sg13g2_FILL8
XSTDFILL110_1056 VDD VSS sg13g2_FILL8
XSTDFILL110_1064 VDD VSS sg13g2_FILL8
XSTDFILL110_1072 VDD VSS sg13g2_FILL8
XSTDFILL110_1080 VDD VSS sg13g2_FILL8
XSTDFILL110_1088 VDD VSS sg13g2_FILL8
XSTDFILL110_1096 VDD VSS sg13g2_FILL8
XSTDFILL110_1104 VDD VSS sg13g2_FILL8
XSTDFILL110_1112 VDD VSS sg13g2_FILL8
XSTDFILL110_1120 VDD VSS sg13g2_FILL8
XSTDFILL110_1128 VDD VSS sg13g2_FILL8
XSTDFILL110_1136 VDD VSS sg13g2_FILL8
XSTDFILL110_1144 VDD VSS sg13g2_FILL8
XSTDFILL110_1152 VDD VSS sg13g2_FILL8
XSTDFILL110_1160 VDD VSS sg13g2_FILL8
XSTDFILL110_1168 VDD VSS sg13g2_FILL8
XSTDFILL110_1176 VDD VSS sg13g2_FILL8
XSTDFILL110_1184 VDD VSS sg13g2_FILL8
XSTDFILL110_1192 VDD VSS sg13g2_FILL8
XSTDFILL110_1200 VDD VSS sg13g2_FILL8
XSTDFILL110_1208 VDD VSS sg13g2_FILL8
XSTDFILL110_1216 VDD VSS sg13g2_FILL8
XSTDFILL110_1224 VDD VSS sg13g2_FILL8
XSTDFILL110_1232 VDD VSS sg13g2_FILL8
XSTDFILL110_1240 VDD VSS sg13g2_FILL8
XSTDFILL110_1248 VDD VSS sg13g2_FILL8
XSTDFILL110_1256 VDD VSS sg13g2_FILL8
XSTDFILL110_1264 VDD VSS sg13g2_FILL8
XSTDFILL110_1272 VDD VSS sg13g2_FILL8
XSTDFILL110_1280 VDD VSS sg13g2_FILL8
XSTDFILL110_1288 VDD VSS sg13g2_FILL8
XSTDFILL110_1296 VDD VSS sg13g2_FILL8
XSTDFILL110_1304 VDD VSS sg13g2_FILL8
XSTDFILL110_1312 VDD VSS sg13g2_FILL8
XSTDFILL110_1320 VDD VSS sg13g2_FILL8
XSTDFILL110_1328 VDD VSS sg13g2_FILL8
XSTDFILL110_1336 VDD VSS sg13g2_FILL8
XSTDFILL110_1344 VDD VSS sg13g2_FILL8
XSTDFILL110_1352 VDD VSS sg13g2_FILL8
XSTDFILL110_1360 VDD VSS sg13g2_FILL8
XSTDFILL110_1368 VDD VSS sg13g2_FILL8
XSTDFILL110_1376 VDD VSS sg13g2_FILL8
XSTDFILL110_1384 VDD VSS sg13g2_FILL8
XSTDFILL110_1392 VDD VSS sg13g2_FILL8
XSTDFILL110_1400 VDD VSS sg13g2_FILL8
XSTDFILL110_1408 VDD VSS sg13g2_FILL8
XSTDFILL110_1416 VDD VSS sg13g2_FILL8
XSTDFILL110_1424 VDD VSS sg13g2_FILL8
XSTDFILL110_1432 VDD VSS sg13g2_FILL8
XSTDFILL110_1440 VDD VSS sg13g2_FILL8
XSTDFILL110_1448 VDD VSS sg13g2_FILL8
XSTDFILL110_1456 VDD VSS sg13g2_FILL8
XSTDFILL110_1464 VDD VSS sg13g2_FILL8
XSTDFILL110_1472 VDD VSS sg13g2_FILL8
XSTDFILL110_1480 VDD VSS sg13g2_FILL8
XSTDFILL110_1488 VDD VSS sg13g2_FILL8
XSTDFILL110_1496 VDD VSS sg13g2_FILL8
XSTDFILL110_1504 VDD VSS sg13g2_FILL8
XSTDFILL110_1512 VDD VSS sg13g2_FILL8
XSTDFILL110_1520 VDD VSS sg13g2_FILL8
XSTDFILL110_1528 VDD VSS sg13g2_FILL2
XSTDFILL110_1530 VDD VSS sg13g2_FILL1
XSTDFILL111_0 VDD VSS sg13g2_FILL8
XSTDFILL111_8 VDD VSS sg13g2_FILL8
XSTDFILL111_16 VDD VSS sg13g2_FILL8
XSTDFILL111_24 VDD VSS sg13g2_FILL8
XSTDFILL111_32 VDD VSS sg13g2_FILL8
XSTDFILL111_40 VDD VSS sg13g2_FILL8
XSTDFILL111_48 VDD VSS sg13g2_FILL8
XSTDFILL111_56 VDD VSS sg13g2_FILL8
XSTDFILL111_64 VDD VSS sg13g2_FILL8
XSTDFILL111_72 VDD VSS sg13g2_FILL8
XSTDFILL111_80 VDD VSS sg13g2_FILL8
XSTDFILL111_88 VDD VSS sg13g2_FILL8
XSTDFILL111_96 VDD VSS sg13g2_FILL8
XSTDFILL111_104 VDD VSS sg13g2_FILL8
XSTDFILL111_112 VDD VSS sg13g2_FILL8
XSTDFILL111_120 VDD VSS sg13g2_FILL8
XSTDFILL111_128 VDD VSS sg13g2_FILL8
XSTDFILL111_136 VDD VSS sg13g2_FILL8
XSTDFILL111_144 VDD VSS sg13g2_FILL8
XSTDFILL111_152 VDD VSS sg13g2_FILL8
XSTDFILL111_160 VDD VSS sg13g2_FILL8
XSTDFILL111_168 VDD VSS sg13g2_FILL8
XSTDFILL111_176 VDD VSS sg13g2_FILL8
XSTDFILL111_184 VDD VSS sg13g2_FILL8
XSTDFILL111_192 VDD VSS sg13g2_FILL8
XSTDFILL111_200 VDD VSS sg13g2_FILL8
XSTDFILL111_208 VDD VSS sg13g2_FILL8
XSTDFILL111_216 VDD VSS sg13g2_FILL8
XSTDFILL111_224 VDD VSS sg13g2_FILL8
XSTDFILL111_232 VDD VSS sg13g2_FILL8
XSTDFILL111_240 VDD VSS sg13g2_FILL8
XSTDFILL111_248 VDD VSS sg13g2_FILL8
XSTDFILL111_256 VDD VSS sg13g2_FILL8
XSTDFILL111_264 VDD VSS sg13g2_FILL8
XSTDFILL111_272 VDD VSS sg13g2_FILL8
XSTDFILL111_280 VDD VSS sg13g2_FILL8
XSTDFILL111_288 VDD VSS sg13g2_FILL8
XSTDFILL111_296 VDD VSS sg13g2_FILL8
XSTDFILL111_304 VDD VSS sg13g2_FILL8
XSTDFILL111_312 VDD VSS sg13g2_FILL8
XSTDFILL111_320 VDD VSS sg13g2_FILL8
XSTDFILL111_328 VDD VSS sg13g2_FILL8
XSTDFILL111_336 VDD VSS sg13g2_FILL8
XSTDFILL111_344 VDD VSS sg13g2_FILL8
XSTDFILL111_352 VDD VSS sg13g2_FILL8
XSTDFILL111_360 VDD VSS sg13g2_FILL8
XSTDFILL111_368 VDD VSS sg13g2_FILL8
XSTDFILL111_376 VDD VSS sg13g2_FILL8
XSTDFILL111_384 VDD VSS sg13g2_FILL8
XSTDFILL111_392 VDD VSS sg13g2_FILL8
XSTDFILL111_400 VDD VSS sg13g2_FILL8
XSTDFILL111_408 VDD VSS sg13g2_FILL8
XSTDFILL111_416 VDD VSS sg13g2_FILL8
XSTDFILL111_424 VDD VSS sg13g2_FILL8
XSTDFILL111_432 VDD VSS sg13g2_FILL8
XSTDFILL111_440 VDD VSS sg13g2_FILL8
XSTDFILL111_448 VDD VSS sg13g2_FILL8
XSTDFILL111_456 VDD VSS sg13g2_FILL8
XSTDFILL111_464 VDD VSS sg13g2_FILL8
XSTDFILL111_472 VDD VSS sg13g2_FILL8
XSTDFILL111_480 VDD VSS sg13g2_FILL8
XSTDFILL111_488 VDD VSS sg13g2_FILL8
XSTDFILL111_496 VDD VSS sg13g2_FILL8
XSTDFILL111_504 VDD VSS sg13g2_FILL8
XSTDFILL111_512 VDD VSS sg13g2_FILL8
XSTDFILL111_520 VDD VSS sg13g2_FILL8
XSTDFILL111_528 VDD VSS sg13g2_FILL8
XSTDFILL111_536 VDD VSS sg13g2_FILL8
XSTDFILL111_544 VDD VSS sg13g2_FILL8
XSTDFILL111_552 VDD VSS sg13g2_FILL8
XSTDFILL111_560 VDD VSS sg13g2_FILL8
XSTDFILL111_568 VDD VSS sg13g2_FILL8
XSTDFILL111_576 VDD VSS sg13g2_FILL8
XSTDFILL111_584 VDD VSS sg13g2_FILL8
XSTDFILL111_592 VDD VSS sg13g2_FILL8
XSTDFILL111_600 VDD VSS sg13g2_FILL8
XSTDFILL111_608 VDD VSS sg13g2_FILL8
XSTDFILL111_616 VDD VSS sg13g2_FILL8
XSTDFILL111_624 VDD VSS sg13g2_FILL8
XSTDFILL111_632 VDD VSS sg13g2_FILL8
XSTDFILL111_640 VDD VSS sg13g2_FILL8
XSTDFILL111_648 VDD VSS sg13g2_FILL8
XSTDFILL111_656 VDD VSS sg13g2_FILL8
XSTDFILL111_664 VDD VSS sg13g2_FILL8
XSTDFILL111_672 VDD VSS sg13g2_FILL8
XSTDFILL111_680 VDD VSS sg13g2_FILL8
XSTDFILL111_688 VDD VSS sg13g2_FILL8
XSTDFILL111_696 VDD VSS sg13g2_FILL8
XSTDFILL111_704 VDD VSS sg13g2_FILL8
XSTDFILL111_712 VDD VSS sg13g2_FILL8
XSTDFILL111_720 VDD VSS sg13g2_FILL8
XSTDFILL111_728 VDD VSS sg13g2_FILL8
XSTDFILL111_736 VDD VSS sg13g2_FILL8
XSTDFILL111_744 VDD VSS sg13g2_FILL8
XSTDFILL111_752 VDD VSS sg13g2_FILL8
XSTDFILL111_760 VDD VSS sg13g2_FILL8
XSTDFILL111_768 VDD VSS sg13g2_FILL8
XSTDFILL111_776 VDD VSS sg13g2_FILL8
XSTDFILL111_784 VDD VSS sg13g2_FILL8
XSTDFILL111_792 VDD VSS sg13g2_FILL8
XSTDFILL111_800 VDD VSS sg13g2_FILL8
XSTDFILL111_808 VDD VSS sg13g2_FILL8
XSTDFILL111_816 VDD VSS sg13g2_FILL8
XSTDFILL111_824 VDD VSS sg13g2_FILL8
XSTDFILL111_832 VDD VSS sg13g2_FILL8
XSTDFILL111_840 VDD VSS sg13g2_FILL8
XSTDFILL111_848 VDD VSS sg13g2_FILL8
XSTDFILL111_856 VDD VSS sg13g2_FILL8
XSTDFILL111_864 VDD VSS sg13g2_FILL8
XSTDFILL111_872 VDD VSS sg13g2_FILL8
XSTDFILL111_880 VDD VSS sg13g2_FILL8
XSTDFILL111_888 VDD VSS sg13g2_FILL8
XSTDFILL111_896 VDD VSS sg13g2_FILL8
XSTDFILL111_904 VDD VSS sg13g2_FILL8
XSTDFILL111_912 VDD VSS sg13g2_FILL8
XSTDFILL111_920 VDD VSS sg13g2_FILL8
XSTDFILL111_928 VDD VSS sg13g2_FILL8
XSTDFILL111_936 VDD VSS sg13g2_FILL8
XSTDFILL111_944 VDD VSS sg13g2_FILL8
XSTDFILL111_952 VDD VSS sg13g2_FILL8
XSTDFILL111_960 VDD VSS sg13g2_FILL8
XSTDFILL111_968 VDD VSS sg13g2_FILL8
XSTDFILL111_976 VDD VSS sg13g2_FILL8
XSTDFILL111_984 VDD VSS sg13g2_FILL8
XSTDFILL111_992 VDD VSS sg13g2_FILL8
XSTDFILL111_1000 VDD VSS sg13g2_FILL8
XSTDFILL111_1008 VDD VSS sg13g2_FILL8
XSTDFILL111_1016 VDD VSS sg13g2_FILL8
XSTDFILL111_1024 VDD VSS sg13g2_FILL8
XSTDFILL111_1032 VDD VSS sg13g2_FILL8
XSTDFILL111_1040 VDD VSS sg13g2_FILL8
XSTDFILL111_1048 VDD VSS sg13g2_FILL8
XSTDFILL111_1056 VDD VSS sg13g2_FILL8
XSTDFILL111_1064 VDD VSS sg13g2_FILL8
XSTDFILL111_1072 VDD VSS sg13g2_FILL8
XSTDFILL111_1080 VDD VSS sg13g2_FILL8
XSTDFILL111_1088 VDD VSS sg13g2_FILL8
XSTDFILL111_1096 VDD VSS sg13g2_FILL8
XSTDFILL111_1104 VDD VSS sg13g2_FILL8
XSTDFILL111_1112 VDD VSS sg13g2_FILL8
XSTDFILL111_1120 VDD VSS sg13g2_FILL8
XSTDFILL111_1128 VDD VSS sg13g2_FILL8
XSTDFILL111_1136 VDD VSS sg13g2_FILL8
XSTDFILL111_1144 VDD VSS sg13g2_FILL8
XSTDFILL111_1152 VDD VSS sg13g2_FILL8
XSTDFILL111_1160 VDD VSS sg13g2_FILL8
XSTDFILL111_1168 VDD VSS sg13g2_FILL8
XSTDFILL111_1176 VDD VSS sg13g2_FILL8
XSTDFILL111_1184 VDD VSS sg13g2_FILL8
XSTDFILL111_1192 VDD VSS sg13g2_FILL8
XSTDFILL111_1200 VDD VSS sg13g2_FILL8
XSTDFILL111_1208 VDD VSS sg13g2_FILL8
XSTDFILL111_1216 VDD VSS sg13g2_FILL8
XSTDFILL111_1224 VDD VSS sg13g2_FILL8
XSTDFILL111_1232 VDD VSS sg13g2_FILL8
XSTDFILL111_1240 VDD VSS sg13g2_FILL8
XSTDFILL111_1248 VDD VSS sg13g2_FILL8
XSTDFILL111_1256 VDD VSS sg13g2_FILL8
XSTDFILL111_1264 VDD VSS sg13g2_FILL8
XSTDFILL111_1272 VDD VSS sg13g2_FILL8
XSTDFILL111_1280 VDD VSS sg13g2_FILL8
XSTDFILL111_1288 VDD VSS sg13g2_FILL8
XSTDFILL111_1296 VDD VSS sg13g2_FILL8
XSTDFILL111_1304 VDD VSS sg13g2_FILL8
XSTDFILL111_1312 VDD VSS sg13g2_FILL8
XSTDFILL111_1320 VDD VSS sg13g2_FILL8
XSTDFILL111_1328 VDD VSS sg13g2_FILL8
XSTDFILL111_1336 VDD VSS sg13g2_FILL8
XSTDFILL111_1344 VDD VSS sg13g2_FILL8
XSTDFILL111_1352 VDD VSS sg13g2_FILL8
XSTDFILL111_1360 VDD VSS sg13g2_FILL8
XSTDFILL111_1368 VDD VSS sg13g2_FILL8
XSTDFILL111_1376 VDD VSS sg13g2_FILL8
XSTDFILL111_1384 VDD VSS sg13g2_FILL8
XSTDFILL111_1392 VDD VSS sg13g2_FILL8
XSTDFILL111_1400 VDD VSS sg13g2_FILL8
XSTDFILL111_1408 VDD VSS sg13g2_FILL8
XSTDFILL111_1416 VDD VSS sg13g2_FILL8
XSTDFILL111_1424 VDD VSS sg13g2_FILL8
XSTDFILL111_1432 VDD VSS sg13g2_FILL8
XSTDFILL111_1440 VDD VSS sg13g2_FILL8
XSTDFILL111_1448 VDD VSS sg13g2_FILL8
XSTDFILL111_1456 VDD VSS sg13g2_FILL8
XSTDFILL111_1464 VDD VSS sg13g2_FILL8
XSTDFILL111_1472 VDD VSS sg13g2_FILL8
XSTDFILL111_1480 VDD VSS sg13g2_FILL8
XSTDFILL111_1488 VDD VSS sg13g2_FILL8
XSTDFILL111_1496 VDD VSS sg13g2_FILL8
XSTDFILL111_1504 VDD VSS sg13g2_FILL8
XSTDFILL111_1512 VDD VSS sg13g2_FILL8
XSTDFILL111_1520 VDD VSS sg13g2_FILL8
XSTDFILL111_1528 VDD VSS sg13g2_FILL2
XSTDFILL111_1530 VDD VSS sg13g2_FILL1
XSTDFILL112_0 VDD VSS sg13g2_FILL8
XSTDFILL112_8 VDD VSS sg13g2_FILL8
XSTDFILL112_16 VDD VSS sg13g2_FILL8
XSTDFILL112_24 VDD VSS sg13g2_FILL8
XSTDFILL112_32 VDD VSS sg13g2_FILL8
XSTDFILL112_40 VDD VSS sg13g2_FILL8
XSTDFILL112_48 VDD VSS sg13g2_FILL8
XSTDFILL112_56 VDD VSS sg13g2_FILL8
XSTDFILL112_64 VDD VSS sg13g2_FILL8
XSTDFILL112_72 VDD VSS sg13g2_FILL8
XSTDFILL112_80 VDD VSS sg13g2_FILL8
XSTDFILL112_88 VDD VSS sg13g2_FILL8
XSTDFILL112_96 VDD VSS sg13g2_FILL8
XSTDFILL112_104 VDD VSS sg13g2_FILL8
XSTDFILL112_112 VDD VSS sg13g2_FILL8
XSTDFILL112_120 VDD VSS sg13g2_FILL8
XSTDFILL112_128 VDD VSS sg13g2_FILL8
XSTDFILL112_136 VDD VSS sg13g2_FILL8
XSTDFILL112_144 VDD VSS sg13g2_FILL8
XSTDFILL112_152 VDD VSS sg13g2_FILL8
XSTDFILL112_160 VDD VSS sg13g2_FILL8
XSTDFILL112_168 VDD VSS sg13g2_FILL8
XSTDFILL112_176 VDD VSS sg13g2_FILL8
XSTDFILL112_184 VDD VSS sg13g2_FILL8
XSTDFILL112_192 VDD VSS sg13g2_FILL8
XSTDFILL112_200 VDD VSS sg13g2_FILL8
XSTDFILL112_208 VDD VSS sg13g2_FILL8
XSTDFILL112_216 VDD VSS sg13g2_FILL8
XSTDFILL112_224 VDD VSS sg13g2_FILL8
XSTDFILL112_232 VDD VSS sg13g2_FILL8
XSTDFILL112_240 VDD VSS sg13g2_FILL8
XSTDFILL112_248 VDD VSS sg13g2_FILL8
XSTDFILL112_256 VDD VSS sg13g2_FILL8
XSTDFILL112_264 VDD VSS sg13g2_FILL8
XSTDFILL112_272 VDD VSS sg13g2_FILL8
XSTDFILL112_280 VDD VSS sg13g2_FILL8
XSTDFILL112_288 VDD VSS sg13g2_FILL8
XSTDFILL112_296 VDD VSS sg13g2_FILL8
XSTDFILL112_304 VDD VSS sg13g2_FILL8
XSTDFILL112_312 VDD VSS sg13g2_FILL8
XSTDFILL112_320 VDD VSS sg13g2_FILL8
XSTDFILL112_328 VDD VSS sg13g2_FILL8
XSTDFILL112_336 VDD VSS sg13g2_FILL8
XSTDFILL112_344 VDD VSS sg13g2_FILL8
XSTDFILL112_352 VDD VSS sg13g2_FILL8
XSTDFILL112_360 VDD VSS sg13g2_FILL8
XSTDFILL112_368 VDD VSS sg13g2_FILL8
XSTDFILL112_376 VDD VSS sg13g2_FILL8
XSTDFILL112_384 VDD VSS sg13g2_FILL8
XSTDFILL112_392 VDD VSS sg13g2_FILL8
XSTDFILL112_400 VDD VSS sg13g2_FILL8
XSTDFILL112_408 VDD VSS sg13g2_FILL8
XSTDFILL112_416 VDD VSS sg13g2_FILL8
XSTDFILL112_424 VDD VSS sg13g2_FILL8
XSTDFILL112_432 VDD VSS sg13g2_FILL8
XSTDFILL112_440 VDD VSS sg13g2_FILL8
XSTDFILL112_448 VDD VSS sg13g2_FILL8
XSTDFILL112_456 VDD VSS sg13g2_FILL8
XSTDFILL112_464 VDD VSS sg13g2_FILL8
XSTDFILL112_472 VDD VSS sg13g2_FILL8
XSTDFILL112_480 VDD VSS sg13g2_FILL8
XSTDFILL112_488 VDD VSS sg13g2_FILL8
XSTDFILL112_496 VDD VSS sg13g2_FILL8
XSTDFILL112_504 VDD VSS sg13g2_FILL8
XSTDFILL112_512 VDD VSS sg13g2_FILL8
XSTDFILL112_520 VDD VSS sg13g2_FILL8
XSTDFILL112_528 VDD VSS sg13g2_FILL8
XSTDFILL112_536 VDD VSS sg13g2_FILL8
XSTDFILL112_544 VDD VSS sg13g2_FILL8
XSTDFILL112_552 VDD VSS sg13g2_FILL8
XSTDFILL112_560 VDD VSS sg13g2_FILL8
XSTDFILL112_568 VDD VSS sg13g2_FILL8
XSTDFILL112_576 VDD VSS sg13g2_FILL8
XSTDFILL112_584 VDD VSS sg13g2_FILL8
XSTDFILL112_592 VDD VSS sg13g2_FILL8
XSTDFILL112_600 VDD VSS sg13g2_FILL8
XSTDFILL112_608 VDD VSS sg13g2_FILL8
XSTDFILL112_616 VDD VSS sg13g2_FILL8
XSTDFILL112_624 VDD VSS sg13g2_FILL8
XSTDFILL112_632 VDD VSS sg13g2_FILL8
XSTDFILL112_640 VDD VSS sg13g2_FILL8
XSTDFILL112_648 VDD VSS sg13g2_FILL8
XSTDFILL112_656 VDD VSS sg13g2_FILL8
XSTDFILL112_664 VDD VSS sg13g2_FILL8
XSTDFILL112_672 VDD VSS sg13g2_FILL8
XSTDFILL112_680 VDD VSS sg13g2_FILL8
XSTDFILL112_688 VDD VSS sg13g2_FILL8
XSTDFILL112_696 VDD VSS sg13g2_FILL8
XSTDFILL112_704 VDD VSS sg13g2_FILL8
XSTDFILL112_712 VDD VSS sg13g2_FILL8
XSTDFILL112_720 VDD VSS sg13g2_FILL8
XSTDFILL112_728 VDD VSS sg13g2_FILL8
XSTDFILL112_736 VDD VSS sg13g2_FILL8
XSTDFILL112_744 VDD VSS sg13g2_FILL8
XSTDFILL112_752 VDD VSS sg13g2_FILL8
XSTDFILL112_760 VDD VSS sg13g2_FILL8
XSTDFILL112_768 VDD VSS sg13g2_FILL8
XSTDFILL112_776 VDD VSS sg13g2_FILL8
XSTDFILL112_784 VDD VSS sg13g2_FILL8
XSTDFILL112_792 VDD VSS sg13g2_FILL8
XSTDFILL112_800 VDD VSS sg13g2_FILL8
XSTDFILL112_808 VDD VSS sg13g2_FILL8
XSTDFILL112_816 VDD VSS sg13g2_FILL8
XSTDFILL112_824 VDD VSS sg13g2_FILL8
XSTDFILL112_832 VDD VSS sg13g2_FILL8
XSTDFILL112_840 VDD VSS sg13g2_FILL8
XSTDFILL112_848 VDD VSS sg13g2_FILL8
XSTDFILL112_856 VDD VSS sg13g2_FILL8
XSTDFILL112_864 VDD VSS sg13g2_FILL8
XSTDFILL112_872 VDD VSS sg13g2_FILL8
XSTDFILL112_880 VDD VSS sg13g2_FILL8
XSTDFILL112_888 VDD VSS sg13g2_FILL8
XSTDFILL112_896 VDD VSS sg13g2_FILL8
XSTDFILL112_904 VDD VSS sg13g2_FILL8
XSTDFILL112_912 VDD VSS sg13g2_FILL8
XSTDFILL112_920 VDD VSS sg13g2_FILL8
XSTDFILL112_928 VDD VSS sg13g2_FILL8
XSTDFILL112_936 VDD VSS sg13g2_FILL8
XSTDFILL112_944 VDD VSS sg13g2_FILL8
XSTDFILL112_952 VDD VSS sg13g2_FILL8
XSTDFILL112_960 VDD VSS sg13g2_FILL8
XSTDFILL112_968 VDD VSS sg13g2_FILL8
XSTDFILL112_976 VDD VSS sg13g2_FILL8
XSTDFILL112_984 VDD VSS sg13g2_FILL8
XSTDFILL112_992 VDD VSS sg13g2_FILL8
XSTDFILL112_1000 VDD VSS sg13g2_FILL8
XSTDFILL112_1008 VDD VSS sg13g2_FILL8
XSTDFILL112_1016 VDD VSS sg13g2_FILL8
XSTDFILL112_1024 VDD VSS sg13g2_FILL8
XSTDFILL112_1032 VDD VSS sg13g2_FILL8
XSTDFILL112_1040 VDD VSS sg13g2_FILL8
XSTDFILL112_1048 VDD VSS sg13g2_FILL8
XSTDFILL112_1056 VDD VSS sg13g2_FILL8
XSTDFILL112_1064 VDD VSS sg13g2_FILL8
XSTDFILL112_1072 VDD VSS sg13g2_FILL8
XSTDFILL112_1080 VDD VSS sg13g2_FILL8
XSTDFILL112_1088 VDD VSS sg13g2_FILL8
XSTDFILL112_1096 VDD VSS sg13g2_FILL8
XSTDFILL112_1104 VDD VSS sg13g2_FILL8
XSTDFILL112_1112 VDD VSS sg13g2_FILL8
XSTDFILL112_1120 VDD VSS sg13g2_FILL8
XSTDFILL112_1128 VDD VSS sg13g2_FILL8
XSTDFILL112_1136 VDD VSS sg13g2_FILL8
XSTDFILL112_1144 VDD VSS sg13g2_FILL8
XSTDFILL112_1152 VDD VSS sg13g2_FILL8
XSTDFILL112_1160 VDD VSS sg13g2_FILL8
XSTDFILL112_1168 VDD VSS sg13g2_FILL8
XSTDFILL112_1176 VDD VSS sg13g2_FILL8
XSTDFILL112_1184 VDD VSS sg13g2_FILL8
XSTDFILL112_1192 VDD VSS sg13g2_FILL8
XSTDFILL112_1200 VDD VSS sg13g2_FILL8
XSTDFILL112_1208 VDD VSS sg13g2_FILL8
XSTDFILL112_1216 VDD VSS sg13g2_FILL8
XSTDFILL112_1224 VDD VSS sg13g2_FILL8
XSTDFILL112_1232 VDD VSS sg13g2_FILL8
XSTDFILL112_1240 VDD VSS sg13g2_FILL8
XSTDFILL112_1248 VDD VSS sg13g2_FILL8
XSTDFILL112_1256 VDD VSS sg13g2_FILL8
XSTDFILL112_1264 VDD VSS sg13g2_FILL8
XSTDFILL112_1272 VDD VSS sg13g2_FILL8
XSTDFILL112_1280 VDD VSS sg13g2_FILL8
XSTDFILL112_1288 VDD VSS sg13g2_FILL8
XSTDFILL112_1296 VDD VSS sg13g2_FILL8
XSTDFILL112_1304 VDD VSS sg13g2_FILL8
XSTDFILL112_1312 VDD VSS sg13g2_FILL8
XSTDFILL112_1320 VDD VSS sg13g2_FILL8
XSTDFILL112_1328 VDD VSS sg13g2_FILL8
XSTDFILL112_1336 VDD VSS sg13g2_FILL8
XSTDFILL112_1344 VDD VSS sg13g2_FILL8
XSTDFILL112_1352 VDD VSS sg13g2_FILL8
XSTDFILL112_1360 VDD VSS sg13g2_FILL8
XSTDFILL112_1368 VDD VSS sg13g2_FILL8
XSTDFILL112_1376 VDD VSS sg13g2_FILL8
XSTDFILL112_1384 VDD VSS sg13g2_FILL8
XSTDFILL112_1392 VDD VSS sg13g2_FILL8
XSTDFILL112_1400 VDD VSS sg13g2_FILL8
XSTDFILL112_1408 VDD VSS sg13g2_FILL8
XSTDFILL112_1416 VDD VSS sg13g2_FILL8
XSTDFILL112_1424 VDD VSS sg13g2_FILL8
XSTDFILL112_1432 VDD VSS sg13g2_FILL8
XSTDFILL112_1440 VDD VSS sg13g2_FILL8
XSTDFILL112_1448 VDD VSS sg13g2_FILL8
XSTDFILL112_1456 VDD VSS sg13g2_FILL8
XSTDFILL112_1464 VDD VSS sg13g2_FILL8
XSTDFILL112_1472 VDD VSS sg13g2_FILL8
XSTDFILL112_1480 VDD VSS sg13g2_FILL8
XSTDFILL112_1488 VDD VSS sg13g2_FILL8
XSTDFILL112_1496 VDD VSS sg13g2_FILL8
XSTDFILL112_1504 VDD VSS sg13g2_FILL8
XSTDFILL112_1512 VDD VSS sg13g2_FILL8
XSTDFILL112_1520 VDD VSS sg13g2_FILL8
XSTDFILL112_1528 VDD VSS sg13g2_FILL2
XSTDFILL112_1530 VDD VSS sg13g2_FILL1
Xseal sealring
.ENDS asicone_202508
