* NGSPICE file created from DCP_DCN_diodes.ext - technology: ihp-sg13g2

.subckt sg13g2_DCNDiode guard anode cathode VSUB
X0 VSUB cathode dantenna l=0 w=0
X1 VSUB cathode dantenna l=0 w=0
C0 cathode anode 3.50574f
C1 guard anode 2.59423f
C2 cathode VSUB 1.7951f
C3 guard VSUB 3.84456f
C4 anode VSUB 8.37275f
.ends

.subckt sg13g2_DCPDiode guard cathode anode
X0 anode cathode dpantenna l=0.16u w=96.87u
X1 anode cathode dpantenna l=0.16u w=96.87u
C0 anode cathode 5.30084f
C1 cathode guard 3.48148f
.ends

.subckt DCP_DCN_diodes VSS VDD guard pad
Xsg13g2_DCNDiode_0 VDD VSS pad VSS sg13g2_DCNDiode
Xsg13g2_DCPDiode_0 VSS VDD pad sg13g2_DCPDiode
C0 VSS pad 0.34356f
C1 VSS guard 5.66987f
C2 VSS VDD 2.92423f
C3 pad guard 10.36676f
C4 pad VDD 0.88307f
C5 VDD guard 8.10709f
C6 VSS 0 9.59075f
C7 guard 0 14.1055f
C8 pad 0 2.38891f
C9 VDD 0 7.35198f
.ends

